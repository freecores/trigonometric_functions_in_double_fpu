
module top_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58;
  wire   [32:0] carry;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  NAND2X1 U1 ( .IN1(n52), .IN2(carry[6]), .QN(n1) );
  NAND2X1 U2 ( .IN1(n57), .IN2(n58), .QN(n2) );
  NAND2X1 U3 ( .IN1(n55), .IN2(carry[3]), .QN(n3) );
  NAND2X1 U4 ( .IN1(B[5]), .IN2(n4), .QN(carry[6]) );
  NAND2X1 U5 ( .IN1(B[2]), .IN2(n2), .QN(carry[3]) );
  NAND2X1 U6 ( .IN1(B[7]), .IN2(n1), .QN(carry[8]) );
  AND2X1 U7 ( .IN1(B[4]), .IN2(n3), .Q(n4) );
  AND2X1 U8 ( .IN1(n50), .IN2(carry[8]), .Q(n5) );
  AND2X1 U9 ( .IN1(n49), .IN2(n5), .Q(n6) );
  AND2X1 U10 ( .IN1(n48), .IN2(n6), .Q(n7) );
  AND2X1 U11 ( .IN1(n47), .IN2(n7), .Q(n8) );
  AND2X1 U12 ( .IN1(n46), .IN2(n8), .Q(n9) );
  AND2X1 U13 ( .IN1(n45), .IN2(n9), .Q(n10) );
  AND2X1 U14 ( .IN1(n44), .IN2(n10), .Q(n11) );
  AND2X1 U15 ( .IN1(n43), .IN2(n11), .Q(n12) );
  AND2X1 U16 ( .IN1(n42), .IN2(n12), .Q(n13) );
  AND2X1 U17 ( .IN1(n41), .IN2(n13), .Q(n14) );
  AND2X1 U18 ( .IN1(n40), .IN2(n14), .Q(n15) );
  AND2X1 U19 ( .IN1(n39), .IN2(n15), .Q(n16) );
  AND2X1 U20 ( .IN1(n38), .IN2(n16), .Q(n17) );
  AND2X1 U21 ( .IN1(n37), .IN2(n17), .Q(n18) );
  AND2X1 U22 ( .IN1(n36), .IN2(n18), .Q(n19) );
  AND2X1 U23 ( .IN1(n35), .IN2(n19), .Q(n20) );
  AND2X1 U24 ( .IN1(n34), .IN2(n20), .Q(n21) );
  AND2X1 U25 ( .IN1(n33), .IN2(n21), .Q(n22) );
  AND2X1 U26 ( .IN1(n32), .IN2(n22), .Q(n23) );
  AND2X1 U27 ( .IN1(n31), .IN2(n23), .Q(n24) );
  AND2X1 U28 ( .IN1(n30), .IN2(n24), .Q(n25) );
  AND2X1 U29 ( .IN1(n29), .IN2(n25), .Q(n26) );
  INVX0 U30 ( .INP(B[1]), .ZN(n57) );
  INVX0 U31 ( .INP(B[3]), .ZN(n55) );
  INVX0 U32 ( .INP(B[6]), .ZN(n52) );
  INVX0 U33 ( .INP(B[8]), .ZN(n50) );
  INVX0 U34 ( .INP(B[9]), .ZN(n49) );
  INVX0 U35 ( .INP(B[10]), .ZN(n48) );
  INVX0 U36 ( .INP(B[11]), .ZN(n47) );
  INVX0 U37 ( .INP(B[12]), .ZN(n46) );
  INVX0 U38 ( .INP(B[13]), .ZN(n45) );
  INVX0 U39 ( .INP(B[14]), .ZN(n44) );
  INVX0 U40 ( .INP(B[15]), .ZN(n43) );
  INVX0 U41 ( .INP(B[16]), .ZN(n42) );
  INVX0 U42 ( .INP(B[17]), .ZN(n41) );
  INVX0 U43 ( .INP(B[18]), .ZN(n40) );
  INVX0 U44 ( .INP(B[19]), .ZN(n39) );
  INVX0 U45 ( .INP(B[20]), .ZN(n38) );
  INVX0 U46 ( .INP(B[21]), .ZN(n37) );
  INVX0 U47 ( .INP(B[22]), .ZN(n36) );
  INVX0 U48 ( .INP(B[23]), .ZN(n35) );
  INVX0 U49 ( .INP(B[24]), .ZN(n34) );
  INVX0 U50 ( .INP(B[25]), .ZN(n33) );
  INVX0 U51 ( .INP(B[26]), .ZN(n32) );
  INVX0 U52 ( .INP(B[27]), .ZN(n31) );
  INVX0 U53 ( .INP(B[28]), .ZN(n30) );
  INVX0 U54 ( .INP(B[29]), .ZN(n29) );
  INVX0 U55 ( .INP(B[30]), .ZN(n28) );
  INVX0 U56 ( .INP(\B[0] ), .ZN(n58) );
  XOR2X1 U57 ( .IN1(B[31]), .IN2(n27), .Q(DIFF[31]) );
  NAND2X1 U58 ( .IN1(n28), .IN2(n26), .QN(n27) );
  INVX0 U59 ( .INP(B[2]), .ZN(n56) );
  INVX0 U60 ( .INP(B[4]), .ZN(n54) );
  INVX0 U61 ( .INP(B[5]), .ZN(n53) );
  INVX0 U62 ( .INP(B[7]), .ZN(n51) );
  XOR2X1 U63 ( .IN1(n1), .IN2(n51), .Q(DIFF[7]) );
  XOR2X1 U64 ( .IN1(n4), .IN2(n53), .Q(DIFF[5]) );
  XOR2X1 U65 ( .IN1(n3), .IN2(n54), .Q(DIFF[4]) );
  XOR2X1 U66 ( .IN1(n2), .IN2(n56), .Q(DIFF[2]) );
  XOR2X1 U67 ( .IN1(n28), .IN2(n26), .Q(DIFF[30]) );
  XOR2X1 U68 ( .IN1(n29), .IN2(n25), .Q(DIFF[29]) );
  XOR2X1 U69 ( .IN1(n30), .IN2(n24), .Q(DIFF[28]) );
  XOR2X1 U70 ( .IN1(n31), .IN2(n23), .Q(DIFF[27]) );
  XOR2X1 U71 ( .IN1(n32), .IN2(n22), .Q(DIFF[26]) );
  XOR2X1 U72 ( .IN1(n33), .IN2(n21), .Q(DIFF[25]) );
  XOR2X1 U73 ( .IN1(n34), .IN2(n20), .Q(DIFF[24]) );
  XOR2X1 U74 ( .IN1(n35), .IN2(n19), .Q(DIFF[23]) );
  XOR2X1 U75 ( .IN1(n36), .IN2(n18), .Q(DIFF[22]) );
  XOR2X1 U76 ( .IN1(n37), .IN2(n17), .Q(DIFF[21]) );
  XOR2X1 U77 ( .IN1(n38), .IN2(n16), .Q(DIFF[20]) );
  XOR2X1 U78 ( .IN1(n39), .IN2(n15), .Q(DIFF[19]) );
  XOR2X1 U79 ( .IN1(n40), .IN2(n14), .Q(DIFF[18]) );
  XOR2X1 U80 ( .IN1(n41), .IN2(n13), .Q(DIFF[17]) );
  XOR2X1 U81 ( .IN1(n42), .IN2(n12), .Q(DIFF[16]) );
  XOR2X1 U82 ( .IN1(n43), .IN2(n11), .Q(DIFF[15]) );
  XOR2X1 U83 ( .IN1(n44), .IN2(n10), .Q(DIFF[14]) );
  XOR2X1 U84 ( .IN1(n45), .IN2(n9), .Q(DIFF[13]) );
  XOR2X1 U85 ( .IN1(n46), .IN2(n8), .Q(DIFF[12]) );
  XOR2X1 U86 ( .IN1(n47), .IN2(n7), .Q(DIFF[11]) );
  XOR2X1 U87 ( .IN1(n48), .IN2(n6), .Q(DIFF[10]) );
  XOR2X1 U88 ( .IN1(n49), .IN2(n5), .Q(DIFF[9]) );
  XOR2X1 U89 ( .IN1(n50), .IN2(carry[8]), .Q(DIFF[8]) );
  XOR2X1 U90 ( .IN1(n52), .IN2(carry[6]), .Q(DIFF[6]) );
  XOR2X1 U91 ( .IN1(n55), .IN2(carry[3]), .Q(DIFF[3]) );
  XOR2X1 U92 ( .IN1(n57), .IN2(n58), .Q(DIFF[1]) );
endmodule


module top_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58;
  wire   [32:0] carry;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  NAND2X1 U1 ( .IN1(n52), .IN2(carry[6]), .QN(n1) );
  NAND2X1 U2 ( .IN1(n55), .IN2(carry[3]), .QN(n2) );
  NAND2X1 U3 ( .IN1(n57), .IN2(n58), .QN(n3) );
  NAND2X1 U4 ( .IN1(B[5]), .IN2(n26), .QN(carry[6]) );
  NAND2X1 U5 ( .IN1(B[2]), .IN2(n3), .QN(carry[3]) );
  NAND2X1 U6 ( .IN1(B[7]), .IN2(n1), .QN(carry[8]) );
  AND2X1 U7 ( .IN1(n50), .IN2(carry[8]), .Q(n4) );
  AND2X1 U8 ( .IN1(n45), .IN2(n9), .Q(n5) );
  AND2X1 U9 ( .IN1(n39), .IN2(n10), .Q(n6) );
  AND2X1 U10 ( .IN1(n33), .IN2(n11), .Q(n7) );
  AND2X1 U11 ( .IN1(n49), .IN2(n4), .Q(n8) );
  AND2X1 U12 ( .IN1(n46), .IN2(n19), .Q(n9) );
  AND2X1 U13 ( .IN1(n40), .IN2(n21), .Q(n10) );
  AND2X1 U14 ( .IN1(n34), .IN2(n23), .Q(n11) );
  AND2X1 U15 ( .IN1(n44), .IN2(n5), .Q(n12) );
  AND2X1 U16 ( .IN1(n38), .IN2(n6), .Q(n13) );
  AND2X1 U17 ( .IN1(n32), .IN2(n7), .Q(n14) );
  AND2X1 U18 ( .IN1(n43), .IN2(n12), .Q(n15) );
  AND2X1 U19 ( .IN1(n37), .IN2(n13), .Q(n16) );
  AND2X1 U20 ( .IN1(n31), .IN2(n14), .Q(n17) );
  AND2X1 U21 ( .IN1(n48), .IN2(n8), .Q(n18) );
  AND2X1 U22 ( .IN1(n47), .IN2(n18), .Q(n19) );
  AND2X1 U23 ( .IN1(n42), .IN2(n15), .Q(n20) );
  AND2X1 U24 ( .IN1(n41), .IN2(n20), .Q(n21) );
  AND2X1 U25 ( .IN1(n36), .IN2(n16), .Q(n22) );
  AND2X1 U26 ( .IN1(n35), .IN2(n22), .Q(n23) );
  AND2X1 U27 ( .IN1(n30), .IN2(n17), .Q(n24) );
  AND2X1 U28 ( .IN1(n29), .IN2(n24), .Q(n25) );
  AND2X1 U29 ( .IN1(B[4]), .IN2(n2), .Q(n26) );
  INVX0 U30 ( .INP(B[3]), .ZN(n55) );
  INVX0 U31 ( .INP(\B[0] ), .ZN(n58) );
  INVX0 U32 ( .INP(B[2]), .ZN(n56) );
  XOR2X1 U33 ( .IN1(B[31]), .IN2(n27), .Q(DIFF[31]) );
  NAND2X1 U34 ( .IN1(n28), .IN2(n25), .QN(n27) );
  INVX0 U35 ( .INP(B[6]), .ZN(n52) );
  INVX0 U36 ( .INP(B[5]), .ZN(n53) );
  INVX0 U37 ( .INP(B[7]), .ZN(n51) );
  INVX0 U38 ( .INP(B[4]), .ZN(n54) );
  INVX0 U39 ( .INP(B[8]), .ZN(n50) );
  INVX0 U40 ( .INP(B[9]), .ZN(n49) );
  INVX0 U41 ( .INP(B[10]), .ZN(n48) );
  INVX0 U42 ( .INP(B[13]), .ZN(n45) );
  INVX0 U43 ( .INP(B[12]), .ZN(n46) );
  INVX0 U44 ( .INP(B[11]), .ZN(n47) );
  INVX0 U45 ( .INP(B[14]), .ZN(n44) );
  INVX0 U46 ( .INP(B[15]), .ZN(n43) );
  INVX0 U47 ( .INP(B[16]), .ZN(n42) );
  INVX0 U48 ( .INP(B[17]), .ZN(n41) );
  INVX0 U49 ( .INP(B[19]), .ZN(n39) );
  INVX0 U50 ( .INP(B[18]), .ZN(n40) );
  INVX0 U51 ( .INP(B[20]), .ZN(n38) );
  INVX0 U52 ( .INP(B[24]), .ZN(n34) );
  INVX0 U53 ( .INP(B[21]), .ZN(n37) );
  INVX0 U54 ( .INP(B[22]), .ZN(n36) );
  INVX0 U55 ( .INP(B[23]), .ZN(n35) );
  INVX0 U56 ( .INP(B[25]), .ZN(n33) );
  INVX0 U57 ( .INP(B[26]), .ZN(n32) );
  INVX0 U58 ( .INP(B[27]), .ZN(n31) );
  INVX0 U59 ( .INP(B[30]), .ZN(n28) );
  INVX0 U60 ( .INP(B[28]), .ZN(n30) );
  INVX0 U61 ( .INP(B[29]), .ZN(n29) );
  XOR2X1 U62 ( .IN1(n1), .IN2(n51), .Q(DIFF[7]) );
  XOR2X1 U63 ( .IN1(n26), .IN2(n53), .Q(DIFF[5]) );
  XOR2X1 U64 ( .IN1(n2), .IN2(n54), .Q(DIFF[4]) );
  XOR2X1 U65 ( .IN1(n3), .IN2(n56), .Q(DIFF[2]) );
  XOR2X1 U66 ( .IN1(n28), .IN2(n25), .Q(DIFF[30]) );
  XOR2X1 U67 ( .IN1(n29), .IN2(n24), .Q(DIFF[29]) );
  XOR2X1 U68 ( .IN1(n30), .IN2(n17), .Q(DIFF[28]) );
  XOR2X1 U69 ( .IN1(n31), .IN2(n14), .Q(DIFF[27]) );
  XOR2X1 U70 ( .IN1(n32), .IN2(n7), .Q(DIFF[26]) );
  XOR2X1 U71 ( .IN1(n33), .IN2(n11), .Q(DIFF[25]) );
  XOR2X1 U72 ( .IN1(n34), .IN2(n23), .Q(DIFF[24]) );
  XOR2X1 U73 ( .IN1(n35), .IN2(n22), .Q(DIFF[23]) );
  XOR2X1 U74 ( .IN1(n36), .IN2(n16), .Q(DIFF[22]) );
  XOR2X1 U75 ( .IN1(n37), .IN2(n13), .Q(DIFF[21]) );
  XOR2X1 U76 ( .IN1(n38), .IN2(n6), .Q(DIFF[20]) );
  XOR2X1 U77 ( .IN1(n39), .IN2(n10), .Q(DIFF[19]) );
  XOR2X1 U78 ( .IN1(n40), .IN2(n21), .Q(DIFF[18]) );
  XOR2X1 U79 ( .IN1(n41), .IN2(n20), .Q(DIFF[17]) );
  XOR2X1 U80 ( .IN1(n42), .IN2(n15), .Q(DIFF[16]) );
  XOR2X1 U81 ( .IN1(n43), .IN2(n12), .Q(DIFF[15]) );
  XOR2X1 U82 ( .IN1(n44), .IN2(n5), .Q(DIFF[14]) );
  XOR2X1 U83 ( .IN1(n45), .IN2(n9), .Q(DIFF[13]) );
  XOR2X1 U84 ( .IN1(n46), .IN2(n19), .Q(DIFF[12]) );
  XOR2X1 U85 ( .IN1(n47), .IN2(n18), .Q(DIFF[11]) );
  XOR2X1 U86 ( .IN1(n48), .IN2(n8), .Q(DIFF[10]) );
  XOR2X1 U87 ( .IN1(n49), .IN2(n4), .Q(DIFF[9]) );
  XOR2X1 U88 ( .IN1(n50), .IN2(carry[8]), .Q(DIFF[8]) );
  XOR2X1 U89 ( .IN1(n52), .IN2(carry[6]), .Q(DIFF[6]) );
  XOR2X1 U90 ( .IN1(n55), .IN2(carry[3]), .Q(DIFF[3]) );
  XOR2X1 U91 ( .IN1(n57), .IN2(n58), .Q(DIFF[1]) );
  INVX0 U92 ( .INP(B[1]), .ZN(n57) );
endmodule


module top_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n48, n49, n50, n51, n52, n53, n54;
  wire   [32:0] carry;
  assign DIFF[1] = A[1];
  assign DIFF[0] = \A[0] ;
  assign \A[0]  = A[0];

  INVX0 U1 ( .INP(carry[30]), .ZN(n45) );
  NAND2X1 U2 ( .IN1(n49), .IN2(n50), .QN(carry[7]) );
  INVX0 U3 ( .INP(n3), .ZN(n49) );
  NAND2X1 U4 ( .IN1(n51), .IN2(n52), .QN(carry[9]) );
  INVX0 U5 ( .INP(n4), .ZN(n51) );
  NAND2X1 U6 ( .IN1(n53), .IN2(n54), .QN(carry[10]) );
  INVX0 U7 ( .INP(carry[9]), .ZN(n53) );
  NAND2X1 U8 ( .IN1(n5), .IN2(n6), .QN(carry[11]) );
  INVX0 U9 ( .INP(carry[10]), .ZN(n5) );
  NAND2X1 U10 ( .IN1(n7), .IN2(n8), .QN(carry[12]) );
  INVX0 U11 ( .INP(carry[11]), .ZN(n7) );
  NAND2X1 U12 ( .IN1(n9), .IN2(n10), .QN(carry[13]) );
  INVX0 U13 ( .INP(carry[12]), .ZN(n9) );
  NAND2X1 U14 ( .IN1(n11), .IN2(n12), .QN(carry[14]) );
  INVX0 U15 ( .INP(carry[13]), .ZN(n11) );
  NAND2X1 U16 ( .IN1(n13), .IN2(n14), .QN(carry[15]) );
  INVX0 U17 ( .INP(carry[14]), .ZN(n13) );
  NAND2X1 U18 ( .IN1(n15), .IN2(n16), .QN(carry[16]) );
  INVX0 U19 ( .INP(carry[15]), .ZN(n15) );
  NAND2X1 U20 ( .IN1(n17), .IN2(n18), .QN(carry[17]) );
  INVX0 U21 ( .INP(carry[16]), .ZN(n17) );
  NAND2X1 U22 ( .IN1(n19), .IN2(n20), .QN(carry[18]) );
  INVX0 U23 ( .INP(carry[17]), .ZN(n19) );
  NAND2X1 U24 ( .IN1(n21), .IN2(n22), .QN(carry[19]) );
  INVX0 U25 ( .INP(carry[18]), .ZN(n21) );
  NAND2X1 U26 ( .IN1(n23), .IN2(n24), .QN(carry[20]) );
  INVX0 U27 ( .INP(carry[19]), .ZN(n23) );
  NAND2X1 U28 ( .IN1(n25), .IN2(n26), .QN(carry[21]) );
  INVX0 U29 ( .INP(carry[20]), .ZN(n25) );
  NAND2X1 U30 ( .IN1(n27), .IN2(n28), .QN(carry[22]) );
  INVX0 U31 ( .INP(carry[21]), .ZN(n27) );
  NAND2X1 U32 ( .IN1(n29), .IN2(n30), .QN(carry[23]) );
  INVX0 U33 ( .INP(carry[22]), .ZN(n29) );
  NAND2X1 U34 ( .IN1(n31), .IN2(n32), .QN(carry[24]) );
  INVX0 U35 ( .INP(carry[23]), .ZN(n31) );
  NAND2X1 U36 ( .IN1(n33), .IN2(n34), .QN(carry[25]) );
  INVX0 U37 ( .INP(carry[24]), .ZN(n33) );
  NAND2X1 U38 ( .IN1(n35), .IN2(n36), .QN(carry[26]) );
  INVX0 U39 ( .INP(carry[25]), .ZN(n35) );
  NAND2X1 U40 ( .IN1(n37), .IN2(n38), .QN(carry[27]) );
  INVX0 U41 ( .INP(carry[26]), .ZN(n37) );
  NAND2X1 U42 ( .IN1(n39), .IN2(n40), .QN(carry[28]) );
  INVX0 U43 ( .INP(carry[27]), .ZN(n39) );
  NAND2X1 U44 ( .IN1(n41), .IN2(n42), .QN(carry[29]) );
  INVX0 U45 ( .INP(carry[28]), .ZN(n41) );
  NAND2X1 U46 ( .IN1(n43), .IN2(n44), .QN(carry[30]) );
  INVX0 U47 ( .INP(carry[29]), .ZN(n43) );
  XOR2X1 U48 ( .IN1(A[31]), .IN2(n1), .Q(DIFF[31]) );
  AND2X1 U49 ( .IN1(n45), .IN2(n46), .Q(n1) );
  AND2X1 U50 ( .IN1(carry[4]), .IN2(A[4]), .Q(n2) );
  NAND2X1 U51 ( .IN1(DIFF[2]), .IN2(n48), .QN(carry[4]) );
  INVX0 U52 ( .INP(A[2]), .ZN(DIFF[2]) );
  INVX0 U53 ( .INP(A[3]), .ZN(n48) );
  INVX0 U54 ( .INP(A[6]), .ZN(n50) );
  INVX0 U55 ( .INP(A[8]), .ZN(n52) );
  INVX0 U56 ( .INP(A[9]), .ZN(n54) );
  INVX0 U57 ( .INP(A[10]), .ZN(n6) );
  INVX0 U58 ( .INP(A[11]), .ZN(n8) );
  INVX0 U59 ( .INP(A[12]), .ZN(n10) );
  INVX0 U60 ( .INP(A[13]), .ZN(n12) );
  INVX0 U61 ( .INP(A[14]), .ZN(n14) );
  INVX0 U62 ( .INP(A[15]), .ZN(n16) );
  INVX0 U63 ( .INP(A[16]), .ZN(n18) );
  INVX0 U64 ( .INP(A[17]), .ZN(n20) );
  INVX0 U65 ( .INP(A[18]), .ZN(n22) );
  INVX0 U66 ( .INP(A[19]), .ZN(n24) );
  INVX0 U67 ( .INP(A[20]), .ZN(n26) );
  INVX0 U68 ( .INP(A[21]), .ZN(n28) );
  INVX0 U69 ( .INP(A[22]), .ZN(n30) );
  INVX0 U70 ( .INP(A[23]), .ZN(n32) );
  INVX0 U71 ( .INP(A[24]), .ZN(n34) );
  INVX0 U72 ( .INP(A[25]), .ZN(n36) );
  INVX0 U73 ( .INP(A[26]), .ZN(n38) );
  INVX0 U74 ( .INP(A[27]), .ZN(n40) );
  INVX0 U75 ( .INP(A[28]), .ZN(n42) );
  INVX0 U76 ( .INP(A[29]), .ZN(n44) );
  INVX0 U77 ( .INP(A[30]), .ZN(n46) );
  AND2X1 U78 ( .IN1(n2), .IN2(A[5]), .Q(n3) );
  AND2X1 U79 ( .IN1(carry[7]), .IN2(A[7]), .Q(n4) );
  XOR2X1 U80 ( .IN1(n6), .IN2(carry[10]), .Q(DIFF[10]) );
  XOR2X1 U81 ( .IN1(n8), .IN2(carry[11]), .Q(DIFF[11]) );
  XOR2X1 U82 ( .IN1(n10), .IN2(carry[12]), .Q(DIFF[12]) );
  XOR2X1 U83 ( .IN1(n12), .IN2(carry[13]), .Q(DIFF[13]) );
  XOR2X1 U84 ( .IN1(n14), .IN2(carry[14]), .Q(DIFF[14]) );
  XOR2X1 U85 ( .IN1(n16), .IN2(carry[15]), .Q(DIFF[15]) );
  XOR2X1 U86 ( .IN1(n18), .IN2(carry[16]), .Q(DIFF[16]) );
  XOR2X1 U87 ( .IN1(n20), .IN2(carry[17]), .Q(DIFF[17]) );
  XOR2X1 U88 ( .IN1(n22), .IN2(carry[18]), .Q(DIFF[18]) );
  XOR2X1 U89 ( .IN1(n24), .IN2(carry[19]), .Q(DIFF[19]) );
  XOR2X1 U90 ( .IN1(n26), .IN2(carry[20]), .Q(DIFF[20]) );
  XOR2X1 U91 ( .IN1(n28), .IN2(carry[21]), .Q(DIFF[21]) );
  XOR2X1 U92 ( .IN1(n30), .IN2(carry[22]), .Q(DIFF[22]) );
  XOR2X1 U93 ( .IN1(n32), .IN2(carry[23]), .Q(DIFF[23]) );
  XOR2X1 U94 ( .IN1(n34), .IN2(carry[24]), .Q(DIFF[24]) );
  XOR2X1 U95 ( .IN1(n36), .IN2(carry[25]), .Q(DIFF[25]) );
  XOR2X1 U96 ( .IN1(n38), .IN2(carry[26]), .Q(DIFF[26]) );
  XOR2X1 U97 ( .IN1(n40), .IN2(carry[27]), .Q(DIFF[27]) );
  XOR2X1 U98 ( .IN1(n42), .IN2(carry[28]), .Q(DIFF[28]) );
  XOR2X1 U99 ( .IN1(n44), .IN2(carry[29]), .Q(DIFF[29]) );
  XOR2X1 U100 ( .IN1(n46), .IN2(carry[30]), .Q(DIFF[30]) );
  XOR2X1 U101 ( .IN1(n48), .IN2(A[2]), .Q(DIFF[3]) );
  XOR2X1 U102 ( .IN1(n50), .IN2(n3), .Q(DIFF[6]) );
  XOR2X1 U103 ( .IN1(n52), .IN2(n4), .Q(DIFF[8]) );
  XOR2X1 U104 ( .IN1(n54), .IN2(carry[9]), .Q(DIFF[9]) );
  XOR2X1 U105 ( .IN1(carry[4]), .IN2(A[4]), .Q(DIFF[4]) );
  XOR2X1 U106 ( .IN1(n2), .IN2(A[5]), .Q(DIFF[5]) );
  XOR2X1 U107 ( .IN1(carry[7]), .IN2(A[7]), .Q(DIFF[7]) );
endmodule


module top_DW01_sub_3 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58;
  wire   [32:0] carry;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  NAND2X1 U1 ( .IN1(n55), .IN2(carry[3]), .QN(n1) );
  NAND2X1 U2 ( .IN1(n57), .IN2(n58), .QN(n2) );
  NAND2X1 U3 ( .IN1(n52), .IN2(carry[6]), .QN(n3) );
  NAND2X1 U4 ( .IN1(B[7]), .IN2(n3), .QN(carry[8]) );
  INVX0 U5 ( .INP(B[3]), .ZN(n55) );
  NAND2X1 U6 ( .IN1(B[5]), .IN2(n26), .QN(carry[6]) );
  NAND2X1 U7 ( .IN1(B[2]), .IN2(n2), .QN(carry[3]) );
  AND2X1 U8 ( .IN1(n50), .IN2(carry[8]), .Q(n4) );
  AND2X1 U9 ( .IN1(n49), .IN2(n4), .Q(n5) );
  AND2X1 U10 ( .IN1(n38), .IN2(n9), .Q(n6) );
  AND2X1 U11 ( .IN1(n34), .IN2(n14), .Q(n7) );
  AND2X1 U12 ( .IN1(n31), .IN2(n11), .Q(n8) );
  AND2X1 U13 ( .IN1(n39), .IN2(n13), .Q(n9) );
  AND2X1 U14 ( .IN1(n33), .IN2(n7), .Q(n10) );
  AND2X1 U15 ( .IN1(n32), .IN2(n10), .Q(n11) );
  AND2X1 U16 ( .IN1(n30), .IN2(n8), .Q(n12) );
  AND2X1 U17 ( .IN1(n40), .IN2(n18), .Q(n13) );
  AND2X1 U18 ( .IN1(n35), .IN2(n16), .Q(n14) );
  AND2X1 U19 ( .IN1(n37), .IN2(n6), .Q(n15) );
  AND2X1 U20 ( .IN1(n36), .IN2(n15), .Q(n16) );
  AND2X1 U21 ( .IN1(n29), .IN2(n12), .Q(n17) );
  AND2X1 U22 ( .IN1(n41), .IN2(n23), .Q(n18) );
  AND2X1 U23 ( .IN1(n46), .IN2(n25), .Q(n19) );
  AND2X1 U24 ( .IN1(n45), .IN2(n19), .Q(n20) );
  AND2X1 U25 ( .IN1(n44), .IN2(n20), .Q(n21) );
  AND2X1 U26 ( .IN1(n43), .IN2(n21), .Q(n22) );
  AND2X1 U27 ( .IN1(n42), .IN2(n22), .Q(n23) );
  AND2X1 U28 ( .IN1(n48), .IN2(n5), .Q(n24) );
  AND2X1 U29 ( .IN1(n47), .IN2(n24), .Q(n25) );
  AND2X1 U30 ( .IN1(B[4]), .IN2(n1), .Q(n26) );
  INVX0 U31 ( .INP(B[7]), .ZN(n51) );
  INVX0 U32 ( .INP(B[2]), .ZN(n56) );
  XOR2X1 U33 ( .IN1(B[31]), .IN2(n27), .Q(DIFF[31]) );
  NAND2X1 U34 ( .IN1(n28), .IN2(n17), .QN(n27) );
  INVX0 U35 ( .INP(B[6]), .ZN(n52) );
  INVX0 U36 ( .INP(B[5]), .ZN(n53) );
  INVX0 U37 ( .INP(B[4]), .ZN(n54) );
  INVX0 U38 ( .INP(B[8]), .ZN(n50) );
  INVX0 U39 ( .INP(B[9]), .ZN(n49) );
  INVX0 U40 ( .INP(B[10]), .ZN(n48) );
  INVX0 U41 ( .INP(B[12]), .ZN(n46) );
  INVX0 U42 ( .INP(B[13]), .ZN(n45) );
  INVX0 U43 ( .INP(B[14]), .ZN(n44) );
  INVX0 U44 ( .INP(B[11]), .ZN(n47) );
  INVX0 U45 ( .INP(B[17]), .ZN(n41) );
  INVX0 U46 ( .INP(B[15]), .ZN(n43) );
  INVX0 U47 ( .INP(B[16]), .ZN(n42) );
  INVX0 U48 ( .INP(B[20]), .ZN(n38) );
  INVX0 U49 ( .INP(B[19]), .ZN(n39) );
  INVX0 U50 ( .INP(B[18]), .ZN(n40) );
  INVX0 U51 ( .INP(B[21]), .ZN(n37) );
  INVX0 U52 ( .INP(B[24]), .ZN(n34) );
  INVX0 U53 ( .INP(B[23]), .ZN(n35) );
  INVX0 U54 ( .INP(B[22]), .ZN(n36) );
  INVX0 U55 ( .INP(B[27]), .ZN(n31) );
  INVX0 U56 ( .INP(B[25]), .ZN(n33) );
  INVX0 U57 ( .INP(B[26]), .ZN(n32) );
  INVX0 U58 ( .INP(B[28]), .ZN(n30) );
  INVX0 U59 ( .INP(B[30]), .ZN(n28) );
  INVX0 U60 ( .INP(B[29]), .ZN(n29) );
  XOR2X1 U61 ( .IN1(n3), .IN2(n51), .Q(DIFF[7]) );
  XOR2X1 U62 ( .IN1(n26), .IN2(n53), .Q(DIFF[5]) );
  XOR2X1 U63 ( .IN1(n1), .IN2(n54), .Q(DIFF[4]) );
  XOR2X1 U64 ( .IN1(n2), .IN2(n56), .Q(DIFF[2]) );
  XOR2X1 U65 ( .IN1(n28), .IN2(n17), .Q(DIFF[30]) );
  XOR2X1 U66 ( .IN1(n29), .IN2(n12), .Q(DIFF[29]) );
  XOR2X1 U67 ( .IN1(n30), .IN2(n8), .Q(DIFF[28]) );
  XOR2X1 U68 ( .IN1(n31), .IN2(n11), .Q(DIFF[27]) );
  XOR2X1 U69 ( .IN1(n32), .IN2(n10), .Q(DIFF[26]) );
  XOR2X1 U70 ( .IN1(n33), .IN2(n7), .Q(DIFF[25]) );
  XOR2X1 U71 ( .IN1(n34), .IN2(n14), .Q(DIFF[24]) );
  XOR2X1 U72 ( .IN1(n35), .IN2(n16), .Q(DIFF[23]) );
  XOR2X1 U73 ( .IN1(n36), .IN2(n15), .Q(DIFF[22]) );
  XOR2X1 U74 ( .IN1(n37), .IN2(n6), .Q(DIFF[21]) );
  XOR2X1 U75 ( .IN1(n38), .IN2(n9), .Q(DIFF[20]) );
  XOR2X1 U76 ( .IN1(n39), .IN2(n13), .Q(DIFF[19]) );
  XOR2X1 U77 ( .IN1(n40), .IN2(n18), .Q(DIFF[18]) );
  XOR2X1 U78 ( .IN1(n41), .IN2(n23), .Q(DIFF[17]) );
  XOR2X1 U79 ( .IN1(n42), .IN2(n22), .Q(DIFF[16]) );
  XOR2X1 U80 ( .IN1(n43), .IN2(n21), .Q(DIFF[15]) );
  XOR2X1 U81 ( .IN1(n44), .IN2(n20), .Q(DIFF[14]) );
  XOR2X1 U82 ( .IN1(n45), .IN2(n19), .Q(DIFF[13]) );
  XOR2X1 U83 ( .IN1(n46), .IN2(n25), .Q(DIFF[12]) );
  XOR2X1 U84 ( .IN1(n47), .IN2(n24), .Q(DIFF[11]) );
  XOR2X1 U85 ( .IN1(n48), .IN2(n5), .Q(DIFF[10]) );
  XOR2X1 U86 ( .IN1(n49), .IN2(n4), .Q(DIFF[9]) );
  XOR2X1 U87 ( .IN1(n50), .IN2(carry[8]), .Q(DIFF[8]) );
  XOR2X1 U88 ( .IN1(n52), .IN2(carry[6]), .Q(DIFF[6]) );
  XOR2X1 U89 ( .IN1(n55), .IN2(carry[3]), .Q(DIFF[3]) );
  XOR2X1 U90 ( .IN1(n57), .IN2(n58), .Q(DIFF[1]) );
  INVX0 U91 ( .INP(\B[0] ), .ZN(n58) );
  INVX0 U92 ( .INP(B[1]), .ZN(n57) );
endmodule


module top_DW01_sub_4 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51;
  wire   [32:0] carry;
  assign DIFF[1] = A[1];
  assign DIFF[0] = \A[0] ;
  assign \A[0]  = A[0];

  FADDX1 U2_3 ( .A(A[3]), .B(1'b1), .CI(A[2]), .CO(carry[4]), .S(DIFF[3]) );
  NAND2X1 U1 ( .IN1(n46), .IN2(n47), .QN(carry[7]) );
  INVX0 U2 ( .INP(n3), .ZN(n46) );
  NAND2X1 U3 ( .IN1(n48), .IN2(n49), .QN(carry[9]) );
  INVX0 U4 ( .INP(n1), .ZN(n48) );
  NAND2X1 U5 ( .IN1(n50), .IN2(n51), .QN(carry[10]) );
  INVX0 U6 ( .INP(carry[9]), .ZN(n50) );
  NAND2X1 U7 ( .IN1(n24), .IN2(n25), .QN(carry[21]) );
  INVX0 U8 ( .INP(carry[20]), .ZN(n24) );
  NAND2X1 U9 ( .IN1(n32), .IN2(n33), .QN(carry[25]) );
  INVX0 U10 ( .INP(carry[24]), .ZN(n32) );
  NAND2X1 U11 ( .IN1(n38), .IN2(n39), .QN(carry[28]) );
  INVX0 U12 ( .INP(carry[27]), .ZN(n38) );
  NAND2X1 U13 ( .IN1(n22), .IN2(n23), .QN(carry[20]) );
  INVX0 U14 ( .INP(carry[19]), .ZN(n22) );
  NAND2X1 U15 ( .IN1(n34), .IN2(n35), .QN(carry[26]) );
  INVX0 U16 ( .INP(carry[25]), .ZN(n34) );
  NAND2X1 U17 ( .IN1(n40), .IN2(n41), .QN(carry[29]) );
  INVX0 U18 ( .INP(carry[28]), .ZN(n40) );
  NAND2X1 U19 ( .IN1(n30), .IN2(n31), .QN(carry[24]) );
  INVX0 U20 ( .INP(carry[23]), .ZN(n30) );
  NAND2X1 U21 ( .IN1(n20), .IN2(n21), .QN(carry[19]) );
  INVX0 U22 ( .INP(carry[18]), .ZN(n20) );
  NAND2X1 U23 ( .IN1(n26), .IN2(n27), .QN(carry[22]) );
  INVX0 U24 ( .INP(carry[21]), .ZN(n26) );
  NAND2X1 U25 ( .IN1(n28), .IN2(n29), .QN(carry[23]) );
  INVX0 U26 ( .INP(carry[22]), .ZN(n28) );
  NAND2X1 U27 ( .IN1(n42), .IN2(n43), .QN(carry[30]) );
  INVX0 U28 ( .INP(carry[29]), .ZN(n42) );
  NAND2X1 U29 ( .IN1(n18), .IN2(n19), .QN(carry[18]) );
  INVX0 U30 ( .INP(carry[17]), .ZN(n18) );
  NAND2X1 U31 ( .IN1(n12), .IN2(n13), .QN(carry[15]) );
  INVX0 U32 ( .INP(carry[14]), .ZN(n12) );
  NAND2X1 U33 ( .IN1(n14), .IN2(n15), .QN(carry[16]) );
  INVX0 U34 ( .INP(carry[15]), .ZN(n14) );
  NAND2X1 U35 ( .IN1(n16), .IN2(n17), .QN(carry[17]) );
  INVX0 U36 ( .INP(carry[16]), .ZN(n16) );
  NAND2X1 U37 ( .IN1(n4), .IN2(n5), .QN(carry[11]) );
  INVX0 U38 ( .INP(carry[10]), .ZN(n4) );
  NAND2X1 U39 ( .IN1(n6), .IN2(n7), .QN(carry[12]) );
  INVX0 U40 ( .INP(carry[11]), .ZN(n6) );
  NAND2X1 U41 ( .IN1(n44), .IN2(n45), .QN(carry[31]) );
  INVX0 U42 ( .INP(carry[30]), .ZN(n44) );
  AND2X1 U43 ( .IN1(carry[7]), .IN2(A[7]), .Q(n1) );
  NAND2X1 U44 ( .IN1(n36), .IN2(n37), .QN(carry[27]) );
  INVX0 U45 ( .INP(carry[26]), .ZN(n36) );
  NAND2X1 U46 ( .IN1(n10), .IN2(n11), .QN(carry[14]) );
  INVX0 U47 ( .INP(carry[13]), .ZN(n10) );
  NAND2X1 U48 ( .IN1(n8), .IN2(n9), .QN(carry[13]) );
  INVX0 U49 ( .INP(carry[12]), .ZN(n8) );
  AND2X1 U50 ( .IN1(carry[4]), .IN2(A[4]), .Q(n2) );
  AND2X1 U51 ( .IN1(n2), .IN2(A[5]), .Q(n3) );
  XNOR2X1 U52 ( .IN1(A[31]), .IN2(carry[31]), .Q(DIFF[31]) );
  INVX0 U53 ( .INP(A[6]), .ZN(n47) );
  INVX0 U54 ( .INP(A[8]), .ZN(n49) );
  INVX0 U55 ( .INP(A[9]), .ZN(n51) );
  INVX0 U56 ( .INP(A[12]), .ZN(n9) );
  INVX0 U57 ( .INP(A[13]), .ZN(n11) );
  INVX0 U58 ( .INP(A[10]), .ZN(n5) );
  INVX0 U59 ( .INP(A[11]), .ZN(n7) );
  INVX0 U60 ( .INP(A[17]), .ZN(n19) );
  INVX0 U61 ( .INP(A[14]), .ZN(n13) );
  INVX0 U62 ( .INP(A[15]), .ZN(n15) );
  INVX0 U63 ( .INP(A[16]), .ZN(n17) );
  INVX0 U64 ( .INP(A[20]), .ZN(n25) );
  INVX0 U65 ( .INP(A[19]), .ZN(n23) );
  INVX0 U66 ( .INP(A[18]), .ZN(n21) );
  INVX0 U67 ( .INP(A[24]), .ZN(n33) );
  INVX0 U68 ( .INP(A[23]), .ZN(n31) );
  INVX0 U69 ( .INP(A[21]), .ZN(n27) );
  INVX0 U70 ( .INP(A[22]), .ZN(n29) );
  INVX0 U71 ( .INP(A[27]), .ZN(n39) );
  INVX0 U72 ( .INP(A[25]), .ZN(n35) );
  INVX0 U73 ( .INP(A[26]), .ZN(n37) );
  INVX0 U74 ( .INP(A[28]), .ZN(n41) );
  INVX0 U75 ( .INP(A[30]), .ZN(n45) );
  INVX0 U76 ( .INP(A[29]), .ZN(n43) );
  INVX0 U77 ( .INP(A[2]), .ZN(DIFF[2]) );
  XOR2X1 U78 ( .IN1(n5), .IN2(carry[10]), .Q(DIFF[10]) );
  XOR2X1 U79 ( .IN1(n7), .IN2(carry[11]), .Q(DIFF[11]) );
  XOR2X1 U80 ( .IN1(n9), .IN2(carry[12]), .Q(DIFF[12]) );
  XOR2X1 U81 ( .IN1(n11), .IN2(carry[13]), .Q(DIFF[13]) );
  XOR2X1 U82 ( .IN1(n13), .IN2(carry[14]), .Q(DIFF[14]) );
  XOR2X1 U83 ( .IN1(n15), .IN2(carry[15]), .Q(DIFF[15]) );
  XOR2X1 U84 ( .IN1(n17), .IN2(carry[16]), .Q(DIFF[16]) );
  XOR2X1 U85 ( .IN1(n19), .IN2(carry[17]), .Q(DIFF[17]) );
  XOR2X1 U86 ( .IN1(n21), .IN2(carry[18]), .Q(DIFF[18]) );
  XOR2X1 U87 ( .IN1(n23), .IN2(carry[19]), .Q(DIFF[19]) );
  XOR2X1 U88 ( .IN1(n25), .IN2(carry[20]), .Q(DIFF[20]) );
  XOR2X1 U89 ( .IN1(n27), .IN2(carry[21]), .Q(DIFF[21]) );
  XOR2X1 U90 ( .IN1(n29), .IN2(carry[22]), .Q(DIFF[22]) );
  XOR2X1 U91 ( .IN1(n31), .IN2(carry[23]), .Q(DIFF[23]) );
  XOR2X1 U92 ( .IN1(n33), .IN2(carry[24]), .Q(DIFF[24]) );
  XOR2X1 U93 ( .IN1(n35), .IN2(carry[25]), .Q(DIFF[25]) );
  XOR2X1 U94 ( .IN1(n37), .IN2(carry[26]), .Q(DIFF[26]) );
  XOR2X1 U95 ( .IN1(n39), .IN2(carry[27]), .Q(DIFF[27]) );
  XOR2X1 U96 ( .IN1(n41), .IN2(carry[28]), .Q(DIFF[28]) );
  XOR2X1 U97 ( .IN1(n43), .IN2(carry[29]), .Q(DIFF[29]) );
  XOR2X1 U98 ( .IN1(n45), .IN2(carry[30]), .Q(DIFF[30]) );
  XOR2X1 U99 ( .IN1(n47), .IN2(n3), .Q(DIFF[6]) );
  XOR2X1 U100 ( .IN1(n49), .IN2(n1), .Q(DIFF[8]) );
  XOR2X1 U101 ( .IN1(n51), .IN2(carry[9]), .Q(DIFF[9]) );
  XOR2X1 U102 ( .IN1(carry[4]), .IN2(A[4]), .Q(DIFF[4]) );
  XOR2X1 U103 ( .IN1(n2), .IN2(A[5]), .Q(DIFF[5]) );
  XOR2X1 U104 ( .IN1(carry[7]), .IN2(A[7]), .Q(DIFF[7]) );
endmodule


module top_DW01_sub_5 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56;
  wire   [32:0] carry;
  assign DIFF[0] = \A[0] ;
  assign \A[0]  = A[0];

  XOR2X1 U1 ( .IN1(n1), .IN2(carry[31]), .Q(DIFF[31]) );
  INVX1 U2 ( .INP(A[31]), .ZN(n1) );
  NAND2X1 U3 ( .IN1(n53), .IN2(n54), .QN(carry[8]) );
  INVX0 U4 ( .INP(carry[7]), .ZN(n53) );
  NAND2X1 U5 ( .IN1(n49), .IN2(n50), .QN(carry[6]) );
  INVX0 U6 ( .INP(carry[5]), .ZN(n49) );
  NAND2X1 U7 ( .IN1(n47), .IN2(n48), .QN(carry[5]) );
  INVX0 U8 ( .INP(n2), .ZN(n47) );
  NAND2X1 U9 ( .IN1(n55), .IN2(n56), .QN(carry[10]) );
  INVX0 U10 ( .INP(n4), .ZN(n55) );
  NAND2X1 U11 ( .IN1(n25), .IN2(n26), .QN(carry[21]) );
  INVX0 U12 ( .INP(carry[20]), .ZN(n25) );
  NAND2X1 U13 ( .IN1(n33), .IN2(n34), .QN(carry[25]) );
  INVX0 U14 ( .INP(carry[24]), .ZN(n33) );
  NAND2X1 U15 ( .IN1(n39), .IN2(n40), .QN(carry[28]) );
  INVX0 U16 ( .INP(carry[27]), .ZN(n39) );
  NAND2X1 U17 ( .IN1(n23), .IN2(n24), .QN(carry[20]) );
  INVX0 U18 ( .INP(carry[19]), .ZN(n23) );
  NAND2X1 U19 ( .IN1(n35), .IN2(n36), .QN(carry[26]) );
  INVX0 U20 ( .INP(carry[25]), .ZN(n35) );
  NAND2X1 U21 ( .IN1(n31), .IN2(n32), .QN(carry[24]) );
  INVX0 U22 ( .INP(carry[23]), .ZN(n31) );
  NAND2X1 U23 ( .IN1(n21), .IN2(n22), .QN(carry[19]) );
  INVX0 U24 ( .INP(carry[18]), .ZN(n21) );
  NAND2X1 U25 ( .IN1(n27), .IN2(n28), .QN(carry[22]) );
  INVX0 U26 ( .INP(carry[21]), .ZN(n27) );
  NAND2X1 U27 ( .IN1(n29), .IN2(n30), .QN(carry[23]) );
  INVX0 U28 ( .INP(carry[22]), .ZN(n29) );
  NAND2X1 U29 ( .IN1(n43), .IN2(n44), .QN(carry[30]) );
  INVX0 U30 ( .INP(carry[29]), .ZN(n43) );
  NAND2X1 U31 ( .IN1(n19), .IN2(n20), .QN(carry[18]) );
  INVX0 U32 ( .INP(carry[17]), .ZN(n19) );
  NAND2X1 U33 ( .IN1(n51), .IN2(n52), .QN(carry[7]) );
  INVX0 U34 ( .INP(carry[6]), .ZN(n51) );
  NAND2X1 U35 ( .IN1(n13), .IN2(n14), .QN(carry[15]) );
  INVX0 U36 ( .INP(carry[14]), .ZN(n13) );
  NAND2X1 U37 ( .IN1(n15), .IN2(n16), .QN(carry[16]) );
  INVX0 U38 ( .INP(carry[15]), .ZN(n15) );
  NAND2X1 U39 ( .IN1(n17), .IN2(n18), .QN(carry[17]) );
  INVX0 U40 ( .INP(carry[16]), .ZN(n17) );
  NAND2X1 U41 ( .IN1(n5), .IN2(n6), .QN(carry[11]) );
  INVX0 U42 ( .INP(carry[10]), .ZN(n5) );
  NAND2X1 U43 ( .IN1(n7), .IN2(n8), .QN(carry[12]) );
  INVX0 U44 ( .INP(carry[11]), .ZN(n7) );
  NAND2X1 U45 ( .IN1(n45), .IN2(n46), .QN(carry[31]) );
  INVX0 U46 ( .INP(carry[30]), .ZN(n45) );
  AND2X1 U47 ( .IN1(n3), .IN2(A[3]), .Q(n2) );
  NAND2X1 U48 ( .IN1(n41), .IN2(n42), .QN(carry[29]) );
  INVX0 U49 ( .INP(carry[28]), .ZN(n41) );
  NAND2X1 U50 ( .IN1(n37), .IN2(n38), .QN(carry[27]) );
  INVX0 U51 ( .INP(carry[26]), .ZN(n37) );
  NAND2X1 U52 ( .IN1(n11), .IN2(n12), .QN(carry[14]) );
  INVX0 U53 ( .INP(carry[13]), .ZN(n11) );
  NAND2X1 U54 ( .IN1(n9), .IN2(n10), .QN(carry[13]) );
  INVX0 U55 ( .INP(carry[12]), .ZN(n9) );
  INVX0 U56 ( .INP(A[7]), .ZN(n54) );
  INVX0 U57 ( .INP(A[1]), .ZN(DIFF[1]) );
  AND2X1 U58 ( .IN1(A[1]), .IN2(A[2]), .Q(n3) );
  AND2X1 U59 ( .IN1(carry[8]), .IN2(A[8]), .Q(n4) );
  INVX0 U60 ( .INP(A[5]), .ZN(n50) );
  INVX0 U61 ( .INP(A[4]), .ZN(n48) );
  INVX0 U62 ( .INP(A[6]), .ZN(n52) );
  INVX0 U63 ( .INP(A[9]), .ZN(n56) );
  INVX0 U64 ( .INP(A[12]), .ZN(n10) );
  INVX0 U65 ( .INP(A[13]), .ZN(n12) );
  INVX0 U66 ( .INP(A[10]), .ZN(n6) );
  INVX0 U67 ( .INP(A[11]), .ZN(n8) );
  INVX0 U68 ( .INP(A[17]), .ZN(n20) );
  INVX0 U69 ( .INP(A[14]), .ZN(n14) );
  INVX0 U70 ( .INP(A[15]), .ZN(n16) );
  INVX0 U71 ( .INP(A[16]), .ZN(n18) );
  INVX0 U72 ( .INP(A[20]), .ZN(n26) );
  INVX0 U73 ( .INP(A[19]), .ZN(n24) );
  INVX0 U74 ( .INP(A[18]), .ZN(n22) );
  INVX0 U75 ( .INP(A[24]), .ZN(n34) );
  INVX0 U76 ( .INP(A[23]), .ZN(n32) );
  INVX0 U77 ( .INP(A[21]), .ZN(n28) );
  INVX0 U78 ( .INP(A[22]), .ZN(n30) );
  INVX0 U79 ( .INP(A[27]), .ZN(n40) );
  INVX0 U80 ( .INP(A[25]), .ZN(n36) );
  INVX0 U81 ( .INP(A[26]), .ZN(n38) );
  INVX0 U82 ( .INP(A[28]), .ZN(n42) );
  INVX0 U83 ( .INP(A[30]), .ZN(n46) );
  INVX0 U84 ( .INP(A[29]), .ZN(n44) );
  XOR2X1 U85 ( .IN1(n6), .IN2(carry[10]), .Q(DIFF[10]) );
  XOR2X1 U86 ( .IN1(n8), .IN2(carry[11]), .Q(DIFF[11]) );
  XOR2X1 U87 ( .IN1(n10), .IN2(carry[12]), .Q(DIFF[12]) );
  XOR2X1 U88 ( .IN1(n12), .IN2(carry[13]), .Q(DIFF[13]) );
  XOR2X1 U89 ( .IN1(n14), .IN2(carry[14]), .Q(DIFF[14]) );
  XOR2X1 U90 ( .IN1(n16), .IN2(carry[15]), .Q(DIFF[15]) );
  XOR2X1 U91 ( .IN1(n18), .IN2(carry[16]), .Q(DIFF[16]) );
  XOR2X1 U92 ( .IN1(n20), .IN2(carry[17]), .Q(DIFF[17]) );
  XOR2X1 U93 ( .IN1(n22), .IN2(carry[18]), .Q(DIFF[18]) );
  XOR2X1 U94 ( .IN1(n24), .IN2(carry[19]), .Q(DIFF[19]) );
  XOR2X1 U95 ( .IN1(n26), .IN2(carry[20]), .Q(DIFF[20]) );
  XOR2X1 U96 ( .IN1(n28), .IN2(carry[21]), .Q(DIFF[21]) );
  XOR2X1 U97 ( .IN1(n30), .IN2(carry[22]), .Q(DIFF[22]) );
  XOR2X1 U98 ( .IN1(n32), .IN2(carry[23]), .Q(DIFF[23]) );
  XOR2X1 U99 ( .IN1(n34), .IN2(carry[24]), .Q(DIFF[24]) );
  XOR2X1 U100 ( .IN1(n36), .IN2(carry[25]), .Q(DIFF[25]) );
  XOR2X1 U101 ( .IN1(n38), .IN2(carry[26]), .Q(DIFF[26]) );
  XOR2X1 U102 ( .IN1(n40), .IN2(carry[27]), .Q(DIFF[27]) );
  XOR2X1 U103 ( .IN1(n42), .IN2(carry[28]), .Q(DIFF[28]) );
  XOR2X1 U104 ( .IN1(n44), .IN2(carry[29]), .Q(DIFF[29]) );
  XOR2X1 U105 ( .IN1(n46), .IN2(carry[30]), .Q(DIFF[30]) );
  XOR2X1 U106 ( .IN1(n48), .IN2(n2), .Q(DIFF[4]) );
  XOR2X1 U107 ( .IN1(n50), .IN2(carry[5]), .Q(DIFF[5]) );
  XOR2X1 U108 ( .IN1(n52), .IN2(carry[6]), .Q(DIFF[6]) );
  XOR2X1 U109 ( .IN1(n54), .IN2(carry[7]), .Q(DIFF[7]) );
  XOR2X1 U110 ( .IN1(n56), .IN2(n4), .Q(DIFF[9]) );
  XOR2X1 U111 ( .IN1(n3), .IN2(A[3]), .Q(DIFF[3]) );
  XOR2X1 U112 ( .IN1(carry[8]), .IN2(A[8]), .Q(DIFF[8]) );
  XOR2X1 U113 ( .IN1(A[1]), .IN2(A[2]), .Q(DIFF[2]) );
endmodule


module top ( enable, degrees, data1, rst, actv, clk );
  input [31:0] degrees;
  output [63:0] data1;
  input [2:0] actv;
  input enable, rst, clk;
  wire   sin_enable, cos_enable, tan_enable, csc_enable, sec_enable,
         cot_enable, N33, N34, N35, N36, N37, N38, N39, N40, N41, N43, N44,
         N50, N51, N52, N54, N55, N60, N61, N62, N63, N64, N65, N66, N67, N68,
         N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82,
         N83, N84, N85, N86, N87, N88, N89, N90, N91, N93, N94, N95, N96, N97,
         N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109,
         N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120,
         N121, N122, N123, N124, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N193, N194, N195, N196, N197, N198, N199, N200,
         N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211,
         N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222,
         N223, N224, N225, N227, N228, N229, N230, N231, N232, N233, N234,
         N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245,
         N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256,
         N257, N258, N292, N293, N294, N295, N296, N297, N298, N299, N300,
         N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311,
         N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322,
         N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333,
         N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344,
         N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355,
         N356, N357, N384, N385, N386, N387, N388, N389, N390, N391, N392,
         N393, N394, N395, N396, N397, N398, N399, N400, N401, N402, N403,
         N404, N405, N406, N407, N408, N409, N410, N411, N412, N413, N414,
         N415, N416, N417, N418, N419, N420, N421, N422, N423, N424, N425,
         N426, N427, N428, N429, N430, N431, N432, N433, N434, N435, N436,
         N437, N438, N439, N440, N441, N442, N443, N444, N445, N446, N447,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n368, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824;
  wire   [1:0] quad;
  wire   [31:0] degrees_tmp2;
  wire   [63:0] data_sin;
  wire   [63:0] data_cos;
  wire   [63:0] data_tan;
  wire   [63:0] data_csc;
  wire   [63:0] data_sec;
  wire   [63:0] data_cot;
  wire   [31:0] divider_out;
  wire   [31:0] degrees_tmp1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;

  DFFX1 tan_enable_reg ( .D(N35), .CLK(clk), .Q(tan_enable) );
  DFFX1 sec_enable_reg ( .D(N37), .CLK(clk), .Q(sec_enable) );
  DFFX1 csc_enable_reg ( .D(N36), .CLK(clk), .Q(csc_enable) );
  DFFX1 cot_enable_reg ( .D(N38), .CLK(clk), .Q(cot_enable) );
  DFFX1 sin_enable_reg ( .D(N33), .CLK(clk), .Q(sin_enable) );
  DFFX1 cos_enable_reg ( .D(N34), .CLK(clk), .Q(cos_enable) );
  DFFX1 \quad_reg[1]  ( .D(N357), .CLK(clk), .Q(quad[1]) );
  DFFX1 \degrees_tmp1_reg[1]  ( .D(n538), .CLK(clk), .Q(n639) );
  DFFX1 \quad_reg[0]  ( .D(N356), .CLK(clk), .Q(quad[0]) );
  DFFX1 \degrees_tmp2_reg[1]  ( .D(N325), .CLK(clk), .Q(degrees_tmp2[1]) );
  DFFX1 \degrees_tmp2_reg[2]  ( .D(N326), .CLK(clk), .Q(degrees_tmp2[2]) );
  DFFX1 \degrees_tmp2_reg[3]  ( .D(N327), .CLK(clk), .Q(degrees_tmp2[3]) );
  DFFX1 \degrees_tmp2_reg[4]  ( .D(N328), .CLK(clk), .Q(degrees_tmp2[4]) );
  DFFX1 \degrees_tmp2_reg[5]  ( .D(N329), .CLK(clk), .Q(degrees_tmp2[5]) );
  DFFX1 \degrees_tmp2_reg[6]  ( .D(N330), .CLK(clk), .Q(degrees_tmp2[6]) );
  DFFX1 \degrees_tmp2_reg[7]  ( .D(N331), .CLK(clk), .Q(degrees_tmp2[7]) );
  DFFX1 \degrees_tmp2_reg[8]  ( .D(N332), .CLK(clk), .Q(degrees_tmp2[8]) );
  DFFX1 \degrees_tmp2_reg[9]  ( .D(N333), .CLK(clk), .Q(degrees_tmp2[9]) );
  DFFX1 \degrees_tmp2_reg[10]  ( .D(N334), .CLK(clk), .Q(degrees_tmp2[10]) );
  DFFX1 \degrees_tmp2_reg[11]  ( .D(N335), .CLK(clk), .Q(degrees_tmp2[11]) );
  DFFX1 \degrees_tmp2_reg[12]  ( .D(N336), .CLK(clk), .Q(degrees_tmp2[12]) );
  DFFX1 \degrees_tmp2_reg[13]  ( .D(N337), .CLK(clk), .Q(degrees_tmp2[13]) );
  DFFX1 \degrees_tmp2_reg[14]  ( .D(N338), .CLK(clk), .Q(degrees_tmp2[14]) );
  DFFX1 \degrees_tmp2_reg[15]  ( .D(N339), .CLK(clk), .Q(degrees_tmp2[15]) );
  DFFX1 \degrees_tmp2_reg[16]  ( .D(N340), .CLK(clk), .Q(degrees_tmp2[16]) );
  DFFX1 \degrees_tmp2_reg[17]  ( .D(N341), .CLK(clk), .Q(degrees_tmp2[17]) );
  DFFX1 \degrees_tmp2_reg[18]  ( .D(N342), .CLK(clk), .Q(degrees_tmp2[18]) );
  DFFX1 \degrees_tmp2_reg[19]  ( .D(N343), .CLK(clk), .Q(degrees_tmp2[19]) );
  DFFX1 \degrees_tmp2_reg[20]  ( .D(N344), .CLK(clk), .Q(degrees_tmp2[20]) );
  DFFX1 \degrees_tmp2_reg[21]  ( .D(N345), .CLK(clk), .Q(degrees_tmp2[21]) );
  DFFX1 \degrees_tmp2_reg[22]  ( .D(N346), .CLK(clk), .Q(degrees_tmp2[22]) );
  DFFX1 \degrees_tmp2_reg[23]  ( .D(N347), .CLK(clk), .Q(degrees_tmp2[23]) );
  DFFX1 \degrees_tmp2_reg[24]  ( .D(N348), .CLK(clk), .Q(degrees_tmp2[24]) );
  DFFX1 \degrees_tmp2_reg[25]  ( .D(N349), .CLK(clk), .Q(degrees_tmp2[25]) );
  DFFX1 \degrees_tmp2_reg[26]  ( .D(N350), .CLK(clk), .Q(degrees_tmp2[26]) );
  DFFX1 \degrees_tmp2_reg[27]  ( .D(N351), .CLK(clk), .Q(degrees_tmp2[27]) );
  DFFX1 \degrees_tmp2_reg[28]  ( .D(N352), .CLK(clk), .Q(degrees_tmp2[28]) );
  DFFX1 \degrees_tmp2_reg[29]  ( .D(N353), .CLK(clk), .Q(degrees_tmp2[29]) );
  DFFX1 \degrees_tmp2_reg[30]  ( .D(N354), .CLK(clk), .Q(degrees_tmp2[30]) );
  DFFX1 \degrees_tmp2_reg[31]  ( .D(N355), .CLK(clk), .Q(degrees_tmp2[31]) );
  DFFX1 \degrees_tmp2_reg[0]  ( .D(N324), .CLK(clk), .Q(degrees_tmp2[0]) );
  DFFX1 \data1_reg[63]  ( .D(N447), .CLK(clk), .Q(data1[63]) );
  DFFX1 \data1_reg[62]  ( .D(N446), .CLK(clk), .Q(data1[62]) );
  DFFX1 \data1_reg[52]  ( .D(N436), .CLK(clk), .Q(data1[52]) );
  DFFX1 \data1_reg[51]  ( .D(N435), .CLK(clk), .Q(data1[51]) );
  DFFX1 \data1_reg[26]  ( .D(N410), .CLK(clk), .Q(data1[26]) );
  DFFX1 \data1_reg[25]  ( .D(N409), .CLK(clk), .Q(data1[25]) );
  DFFX1 \data1_reg[24]  ( .D(N408), .CLK(clk), .Q(data1[24]) );
  DFFX1 \data1_reg[23]  ( .D(N407), .CLK(clk), .Q(data1[23]) );
  DFFX1 \data1_reg[22]  ( .D(N406), .CLK(clk), .Q(data1[22]) );
  DFFX1 \data1_reg[21]  ( .D(N405), .CLK(clk), .Q(data1[21]) );
  DFFX1 \data1_reg[20]  ( .D(N404), .CLK(clk), .Q(data1[20]) );
  DFFX1 \data1_reg[19]  ( .D(N403), .CLK(clk), .Q(data1[19]) );
  DFFX1 \data1_reg[18]  ( .D(N402), .CLK(clk), .Q(data1[18]) );
  DFFX1 \data1_reg[17]  ( .D(N401), .CLK(clk), .Q(data1[17]) );
  DFFX1 \data1_reg[16]  ( .D(N400), .CLK(clk), .Q(data1[16]) );
  DFFX1 \data1_reg[15]  ( .D(N399), .CLK(clk), .Q(data1[15]) );
  DFFX1 \data1_reg[14]  ( .D(N398), .CLK(clk), .Q(data1[14]) );
  DFFX1 \data1_reg[13]  ( .D(N397), .CLK(clk), .Q(data1[13]) );
  DFFX1 \data1_reg[12]  ( .D(N396), .CLK(clk), .Q(data1[12]) );
  DFFX1 \data1_reg[11]  ( .D(N395), .CLK(clk), .Q(data1[11]) );
  DFFX1 \data1_reg[10]  ( .D(N394), .CLK(clk), .Q(data1[10]) );
  DFFX1 \data1_reg[9]  ( .D(N393), .CLK(clk), .Q(data1[9]) );
  DFFX1 \data1_reg[8]  ( .D(N392), .CLK(clk), .Q(data1[8]) );
  DFFX1 \data1_reg[7]  ( .D(N391), .CLK(clk), .Q(data1[7]) );
  DFFX1 \data1_reg[6]  ( .D(N390), .CLK(clk), .Q(data1[6]) );
  DFFX1 \data1_reg[5]  ( .D(N389), .CLK(clk), .Q(data1[5]) );
  DFFX1 \data1_reg[4]  ( .D(N388), .CLK(clk), .Q(data1[4]) );
  DFFX1 \data1_reg[3]  ( .D(N387), .CLK(clk), .Q(data1[3]) );
  DFFX1 \data1_reg[2]  ( .D(N386), .CLK(clk), .Q(data1[2]) );
  DFFX1 \data1_reg[1]  ( .D(N385), .CLK(clk), .Q(data1[1]) );
  DFFX1 \data1_reg[0]  ( .D(N384), .CLK(clk), .Q(data1[0]) );
  AO22X1 U149 ( .IN1(N193), .IN2(n678), .IN3(degrees_tmp1[0]), .IN4(n679), .Q(
        n537) );
  AO22X1 U151 ( .IN1(N195), .IN2(n678), .IN3(degrees_tmp1[2]), .IN4(n679), .Q(
        n539) );
  AO22X1 U152 ( .IN1(N196), .IN2(n678), .IN3(degrees_tmp1[3]), .IN4(n679), .Q(
        n540) );
  AO22X1 U153 ( .IN1(N197), .IN2(n678), .IN3(degrees_tmp1[4]), .IN4(n679), .Q(
        n541) );
  AO22X1 U154 ( .IN1(N198), .IN2(n678), .IN3(degrees_tmp1[5]), .IN4(n679), .Q(
        n542) );
  AO22X1 U155 ( .IN1(N199), .IN2(n678), .IN3(degrees_tmp1[6]), .IN4(n679), .Q(
        n543) );
  AO22X1 U156 ( .IN1(N200), .IN2(n678), .IN3(degrees_tmp1[7]), .IN4(n679), .Q(
        n544) );
  AO22X1 U157 ( .IN1(N201), .IN2(n678), .IN3(degrees_tmp1[8]), .IN4(n679), .Q(
        n545) );
  AO22X1 U158 ( .IN1(N202), .IN2(n678), .IN3(degrees_tmp1[9]), .IN4(n679), .Q(
        n546) );
  AO22X1 U159 ( .IN1(N203), .IN2(n678), .IN3(degrees_tmp1[10]), .IN4(n679), 
        .Q(n547) );
  AO22X1 U160 ( .IN1(N204), .IN2(n678), .IN3(degrees_tmp1[11]), .IN4(n679), 
        .Q(n548) );
  AO22X1 U161 ( .IN1(N205), .IN2(n678), .IN3(degrees_tmp1[12]), .IN4(n679), 
        .Q(n549) );
  AO22X1 U162 ( .IN1(N206), .IN2(n678), .IN3(degrees_tmp1[13]), .IN4(n679), 
        .Q(n550) );
  AO22X1 U163 ( .IN1(N207), .IN2(n678), .IN3(degrees_tmp1[14]), .IN4(n679), 
        .Q(n551) );
  AO22X1 U164 ( .IN1(N208), .IN2(n224), .IN3(degrees_tmp1[15]), .IN4(n679), 
        .Q(n552) );
  AO22X1 U165 ( .IN1(N209), .IN2(n224), .IN3(degrees_tmp1[16]), .IN4(n679), 
        .Q(n553) );
  AO22X1 U166 ( .IN1(N210), .IN2(n224), .IN3(degrees_tmp1[17]), .IN4(n679), 
        .Q(n554) );
  AO22X1 U167 ( .IN1(N211), .IN2(n224), .IN3(degrees_tmp1[18]), .IN4(n679), 
        .Q(n555) );
  AO22X1 U168 ( .IN1(N212), .IN2(n224), .IN3(degrees_tmp1[19]), .IN4(n679), 
        .Q(n556) );
  AO22X1 U169 ( .IN1(N213), .IN2(n224), .IN3(degrees_tmp1[20]), .IN4(n679), 
        .Q(n557) );
  AO22X1 U170 ( .IN1(N214), .IN2(n224), .IN3(degrees_tmp1[21]), .IN4(n679), 
        .Q(n558) );
  AO22X1 U171 ( .IN1(N215), .IN2(n224), .IN3(degrees_tmp1[22]), .IN4(n679), 
        .Q(n559) );
  AO22X1 U172 ( .IN1(N216), .IN2(n678), .IN3(degrees_tmp1[23]), .IN4(n679), 
        .Q(n560) );
  AO22X1 U173 ( .IN1(N217), .IN2(n224), .IN3(degrees_tmp1[24]), .IN4(n679), 
        .Q(n561) );
  AO22X1 U174 ( .IN1(N218), .IN2(n678), .IN3(degrees_tmp1[25]), .IN4(n679), 
        .Q(n562) );
  AO22X1 U175 ( .IN1(N219), .IN2(n224), .IN3(degrees_tmp1[26]), .IN4(n679), 
        .Q(n563) );
  AO22X1 U176 ( .IN1(N220), .IN2(n224), .IN3(degrees_tmp1[27]), .IN4(n679), 
        .Q(n564) );
  AO22X1 U177 ( .IN1(N221), .IN2(n678), .IN3(degrees_tmp1[28]), .IN4(n679), 
        .Q(n565) );
  AO22X1 U178 ( .IN1(N222), .IN2(n224), .IN3(degrees_tmp1[29]), .IN4(n679), 
        .Q(n566) );
  AO22X1 U179 ( .IN1(N223), .IN2(n678), .IN3(degrees_tmp1[30]), .IN4(n679), 
        .Q(n567) );
  AO22X1 U180 ( .IN1(N224), .IN2(n224), .IN3(degrees_tmp1[31]), .IN4(n679), 
        .Q(n568) );
  AOI222X1 U181 ( .IN1(data_csc[63]), .IN2(n821), .IN3(data_cot[63]), .IN4(
        n654), .IN5(data_sec[63]), .IN6(n658), .QN(n226) );
  AOI222X1 U182 ( .IN1(data_sin[63]), .IN2(n820), .IN3(data_tan[63]), .IN4(
        n649), .IN5(data_cos[63]), .IN6(n645), .QN(n225) );
  AOI222X1 U183 ( .IN1(data_csc[62]), .IN2(n821), .IN3(data_cot[62]), .IN4(
        n655), .IN5(data_sec[62]), .IN6(n659), .QN(n228) );
  AOI222X1 U185 ( .IN1(data_csc[61]), .IN2(n821), .IN3(data_cot[61]), .IN4(
        n656), .IN5(data_sec[61]), .IN6(n660), .QN(n230) );
  AOI222X1 U186 ( .IN1(data_sin[61]), .IN2(n820), .IN3(data_tan[61]), .IN4(
        n649), .IN5(data_cos[61]), .IN6(n646), .QN(n229) );
  AOI222X1 U187 ( .IN1(data_csc[60]), .IN2(n821), .IN3(data_cot[60]), .IN4(
        n657), .IN5(data_sec[60]), .IN6(n661), .QN(n232) );
  AOI222X1 U188 ( .IN1(data_sin[60]), .IN2(n820), .IN3(data_tan[60]), .IN4(
        n649), .IN5(data_cos[60]), .IN6(n647), .QN(n231) );
  AOI222X1 U189 ( .IN1(data_csc[59]), .IN2(n821), .IN3(data_cot[59]), .IN4(
        n657), .IN5(data_sec[59]), .IN6(n658), .QN(n234) );
  AOI222X1 U190 ( .IN1(data_sin[59]), .IN2(n820), .IN3(data_tan[59]), .IN4(
        n649), .IN5(data_cos[59]), .IN6(n648), .QN(n233) );
  AOI222X1 U191 ( .IN1(data_csc[58]), .IN2(n821), .IN3(data_cot[58]), .IN4(
        n657), .IN5(data_sec[58]), .IN6(n659), .QN(n236) );
  AOI222X1 U192 ( .IN1(data_sin[58]), .IN2(n820), .IN3(data_tan[58]), .IN4(
        n649), .IN5(data_cos[58]), .IN6(n648), .QN(n235) );
  AOI222X1 U193 ( .IN1(data_csc[57]), .IN2(n821), .IN3(data_cot[57]), .IN4(
        n657), .IN5(data_sec[57]), .IN6(n660), .QN(n238) );
  AOI222X1 U194 ( .IN1(data_sin[57]), .IN2(n820), .IN3(data_tan[57]), .IN4(
        n649), .IN5(data_cos[57]), .IN6(n648), .QN(n237) );
  AOI222X1 U195 ( .IN1(data_csc[56]), .IN2(n821), .IN3(data_cot[56]), .IN4(
        n657), .IN5(data_sec[56]), .IN6(n661), .QN(n240) );
  AOI222X1 U196 ( .IN1(data_sin[56]), .IN2(n820), .IN3(data_tan[56]), .IN4(
        n649), .IN5(data_cos[56]), .IN6(n648), .QN(n239) );
  AOI222X1 U197 ( .IN1(data_csc[55]), .IN2(n821), .IN3(data_cot[55]), .IN4(
        n657), .IN5(data_sec[55]), .IN6(n658), .QN(n242) );
  AOI222X1 U198 ( .IN1(data_sin[55]), .IN2(n820), .IN3(data_tan[55]), .IN4(
        n649), .IN5(data_cos[55]), .IN6(n648), .QN(n241) );
  AOI222X1 U199 ( .IN1(data_csc[54]), .IN2(n821), .IN3(data_cot[54]), .IN4(
        n657), .IN5(data_sec[54]), .IN6(n659), .QN(n244) );
  AOI222X1 U200 ( .IN1(data_sin[54]), .IN2(n820), .IN3(data_tan[54]), .IN4(
        n649), .IN5(data_cos[54]), .IN6(n648), .QN(n243) );
  AOI222X1 U201 ( .IN1(data_csc[53]), .IN2(n821), .IN3(data_cot[53]), .IN4(
        n657), .IN5(data_sec[53]), .IN6(n660), .QN(n246) );
  AOI222X1 U202 ( .IN1(data_sin[53]), .IN2(n820), .IN3(data_tan[53]), .IN4(
        n649), .IN5(data_cos[53]), .IN6(n648), .QN(n245) );
  AOI222X1 U203 ( .IN1(data_csc[52]), .IN2(n821), .IN3(data_cot[52]), .IN4(
        n657), .IN5(data_sec[52]), .IN6(n661), .QN(n248) );
  AOI222X1 U204 ( .IN1(data_sin[52]), .IN2(n820), .IN3(data_tan[52]), .IN4(
        n649), .IN5(data_cos[52]), .IN6(n648), .QN(n247) );
  AOI222X1 U205 ( .IN1(data_csc[51]), .IN2(n651), .IN3(data_cot[51]), .IN4(
        n657), .IN5(data_sec[51]), .IN6(n658), .QN(n250) );
  AOI222X1 U206 ( .IN1(data_sin[51]), .IN2(n820), .IN3(data_tan[51]), .IN4(
        n649), .IN5(data_cos[51]), .IN6(n648), .QN(n249) );
  AOI222X1 U207 ( .IN1(data_csc[50]), .IN2(n652), .IN3(data_cot[50]), .IN4(
        n657), .IN5(data_sec[50]), .IN6(n659), .QN(n252) );
  AOI222X1 U208 ( .IN1(data_sin[50]), .IN2(n642), .IN3(data_tan[50]), .IN4(
        n649), .IN5(data_cos[50]), .IN6(n648), .QN(n251) );
  AOI222X1 U209 ( .IN1(data_csc[49]), .IN2(n653), .IN3(data_cot[49]), .IN4(
        n657), .IN5(data_sec[49]), .IN6(n660), .QN(n254) );
  AOI222X1 U210 ( .IN1(data_sin[49]), .IN2(n643), .IN3(data_tan[49]), .IN4(
        n649), .IN5(data_cos[49]), .IN6(n648), .QN(n253) );
  AOI222X1 U211 ( .IN1(data_csc[48]), .IN2(n821), .IN3(data_cot[48]), .IN4(
        n657), .IN5(data_sec[48]), .IN6(n661), .QN(n256) );
  AOI222X1 U212 ( .IN1(data_sin[48]), .IN2(n644), .IN3(data_tan[48]), .IN4(
        n649), .IN5(data_cos[48]), .IN6(n648), .QN(n255) );
  AOI222X1 U213 ( .IN1(data_csc[47]), .IN2(n651), .IN3(data_cot[47]), .IN4(
        n654), .IN5(data_sec[47]), .IN6(n661), .QN(n258) );
  AOI222X1 U214 ( .IN1(data_sin[47]), .IN2(n820), .IN3(data_tan[47]), .IN4(
        n649), .IN5(data_cos[47]), .IN6(n648), .QN(n257) );
  AOI222X1 U215 ( .IN1(data_csc[46]), .IN2(n652), .IN3(data_cot[46]), .IN4(
        n655), .IN5(data_sec[46]), .IN6(n661), .QN(n260) );
  AOI222X1 U216 ( .IN1(data_sin[46]), .IN2(n642), .IN3(data_tan[46]), .IN4(
        n649), .IN5(data_cos[46]), .IN6(n645), .QN(n259) );
  AOI222X1 U217 ( .IN1(data_csc[45]), .IN2(n653), .IN3(data_cot[45]), .IN4(
        n656), .IN5(data_sec[45]), .IN6(n661), .QN(n262) );
  AOI222X1 U218 ( .IN1(data_sin[45]), .IN2(n643), .IN3(data_tan[45]), .IN4(
        n649), .IN5(data_cos[45]), .IN6(n646), .QN(n261) );
  AOI222X1 U219 ( .IN1(data_csc[44]), .IN2(n821), .IN3(data_cot[44]), .IN4(
        n657), .IN5(data_sec[44]), .IN6(n661), .QN(n264) );
  AOI222X1 U220 ( .IN1(data_sin[44]), .IN2(n644), .IN3(data_tan[44]), .IN4(
        n649), .IN5(data_cos[44]), .IN6(n647), .QN(n263) );
  AOI222X1 U221 ( .IN1(data_csc[43]), .IN2(n651), .IN3(data_cot[43]), .IN4(
        n654), .IN5(data_sec[43]), .IN6(n661), .QN(n266) );
  AOI222X1 U222 ( .IN1(data_sin[43]), .IN2(n820), .IN3(data_tan[43]), .IN4(
        n649), .IN5(data_cos[43]), .IN6(n648), .QN(n265) );
  AOI222X1 U223 ( .IN1(data_csc[42]), .IN2(n652), .IN3(data_cot[42]), .IN4(
        n655), .IN5(data_sec[42]), .IN6(n661), .QN(n268) );
  AOI222X1 U224 ( .IN1(data_sin[42]), .IN2(n642), .IN3(data_tan[42]), .IN4(
        n649), .IN5(data_cos[42]), .IN6(n645), .QN(n267) );
  AOI222X1 U225 ( .IN1(data_csc[41]), .IN2(n653), .IN3(data_cot[41]), .IN4(
        n656), .IN5(data_sec[41]), .IN6(n661), .QN(n270) );
  AOI222X1 U226 ( .IN1(data_sin[41]), .IN2(n643), .IN3(data_tan[41]), .IN4(
        n649), .IN5(data_cos[41]), .IN6(n646), .QN(n269) );
  AOI222X1 U227 ( .IN1(data_csc[40]), .IN2(n821), .IN3(data_cot[40]), .IN4(
        n657), .IN5(data_sec[40]), .IN6(n661), .QN(n272) );
  AOI222X1 U228 ( .IN1(data_sin[40]), .IN2(n644), .IN3(data_tan[40]), .IN4(
        n649), .IN5(data_cos[40]), .IN6(n647), .QN(n271) );
  AOI222X1 U229 ( .IN1(data_csc[39]), .IN2(n651), .IN3(data_cot[39]), .IN4(
        n654), .IN5(data_sec[39]), .IN6(n661), .QN(n274) );
  AOI222X1 U230 ( .IN1(data_sin[39]), .IN2(n820), .IN3(data_tan[39]), .IN4(
        n649), .IN5(data_cos[39]), .IN6(n648), .QN(n273) );
  AOI222X1 U231 ( .IN1(data_csc[38]), .IN2(n652), .IN3(data_cot[38]), .IN4(
        n655), .IN5(data_sec[38]), .IN6(n661), .QN(n276) );
  AOI222X1 U232 ( .IN1(data_sin[38]), .IN2(n642), .IN3(data_tan[38]), .IN4(
        n649), .IN5(data_cos[38]), .IN6(n645), .QN(n275) );
  AOI222X1 U233 ( .IN1(data_csc[37]), .IN2(n653), .IN3(data_cot[37]), .IN4(
        n656), .IN5(data_sec[37]), .IN6(n661), .QN(n278) );
  AOI222X1 U234 ( .IN1(data_sin[37]), .IN2(n643), .IN3(data_tan[37]), .IN4(
        n649), .IN5(data_cos[37]), .IN6(n646), .QN(n277) );
  AOI222X1 U235 ( .IN1(data_csc[36]), .IN2(n821), .IN3(data_cot[36]), .IN4(
        n657), .IN5(data_sec[36]), .IN6(n661), .QN(n280) );
  AOI222X1 U236 ( .IN1(data_sin[36]), .IN2(n644), .IN3(data_tan[36]), .IN4(
        n649), .IN5(data_cos[36]), .IN6(n647), .QN(n279) );
  AOI222X1 U237 ( .IN1(data_csc[35]), .IN2(n653), .IN3(data_cot[35]), .IN4(
        n656), .IN5(data_sec[35]), .IN6(n660), .QN(n282) );
  AOI222X1 U238 ( .IN1(data_sin[35]), .IN2(n644), .IN3(data_tan[35]), .IN4(
        n649), .IN5(data_cos[35]), .IN6(n647), .QN(n281) );
  AOI222X1 U239 ( .IN1(data_csc[34]), .IN2(n653), .IN3(data_cot[34]), .IN4(
        n656), .IN5(data_sec[34]), .IN6(n660), .QN(n284) );
  AOI222X1 U240 ( .IN1(data_sin[34]), .IN2(n644), .IN3(data_tan[34]), .IN4(
        n649), .IN5(data_cos[34]), .IN6(n647), .QN(n283) );
  AOI222X1 U241 ( .IN1(data_csc[33]), .IN2(n653), .IN3(data_cot[33]), .IN4(
        n656), .IN5(data_sec[33]), .IN6(n660), .QN(n286) );
  AOI222X1 U242 ( .IN1(data_sin[33]), .IN2(n644), .IN3(data_tan[33]), .IN4(
        n649), .IN5(data_cos[33]), .IN6(n647), .QN(n285) );
  AOI222X1 U243 ( .IN1(data_csc[32]), .IN2(n653), .IN3(data_cot[32]), .IN4(
        n656), .IN5(data_sec[32]), .IN6(n660), .QN(n288) );
  AOI222X1 U244 ( .IN1(data_sin[32]), .IN2(n644), .IN3(data_tan[32]), .IN4(
        n649), .IN5(data_cos[32]), .IN6(n647), .QN(n287) );
  AOI222X1 U245 ( .IN1(data_csc[31]), .IN2(n653), .IN3(data_cot[31]), .IN4(
        n656), .IN5(data_sec[31]), .IN6(n660), .QN(n290) );
  AOI222X1 U246 ( .IN1(data_sin[31]), .IN2(n644), .IN3(data_tan[31]), .IN4(
        n649), .IN5(data_cos[31]), .IN6(n647), .QN(n289) );
  AOI222X1 U247 ( .IN1(data_csc[30]), .IN2(n653), .IN3(data_cot[30]), .IN4(
        n656), .IN5(data_sec[30]), .IN6(n660), .QN(n292) );
  AOI222X1 U248 ( .IN1(data_sin[30]), .IN2(n644), .IN3(data_tan[30]), .IN4(
        n649), .IN5(data_cos[30]), .IN6(n647), .QN(n291) );
  AOI222X1 U249 ( .IN1(data_csc[29]), .IN2(n653), .IN3(data_cot[29]), .IN4(
        n656), .IN5(data_sec[29]), .IN6(n660), .QN(n294) );
  AOI222X1 U250 ( .IN1(data_sin[29]), .IN2(n644), .IN3(data_tan[29]), .IN4(
        n650), .IN5(data_cos[29]), .IN6(n647), .QN(n293) );
  AOI222X1 U251 ( .IN1(data_csc[28]), .IN2(n653), .IN3(data_cot[28]), .IN4(
        n656), .IN5(data_sec[28]), .IN6(n660), .QN(n296) );
  AOI222X1 U252 ( .IN1(data_sin[28]), .IN2(n644), .IN3(data_tan[28]), .IN4(
        n650), .IN5(data_cos[28]), .IN6(n647), .QN(n295) );
  AOI222X1 U253 ( .IN1(data_csc[27]), .IN2(n653), .IN3(data_cot[27]), .IN4(
        n656), .IN5(data_sec[27]), .IN6(n660), .QN(n298) );
  AOI222X1 U254 ( .IN1(data_sin[27]), .IN2(n644), .IN3(data_tan[27]), .IN4(
        n650), .IN5(data_cos[27]), .IN6(n647), .QN(n297) );
  AOI222X1 U255 ( .IN1(data_csc[26]), .IN2(n653), .IN3(data_cot[26]), .IN4(
        n656), .IN5(data_sec[26]), .IN6(n660), .QN(n300) );
  AOI222X1 U256 ( .IN1(data_sin[26]), .IN2(n644), .IN3(data_tan[26]), .IN4(
        n650), .IN5(data_cos[26]), .IN6(n647), .QN(n299) );
  AOI222X1 U257 ( .IN1(data_csc[25]), .IN2(n653), .IN3(data_cot[25]), .IN4(
        n656), .IN5(data_sec[25]), .IN6(n660), .QN(n302) );
  AOI222X1 U258 ( .IN1(data_sin[25]), .IN2(n644), .IN3(data_tan[25]), .IN4(
        n650), .IN5(data_cos[25]), .IN6(n647), .QN(n301) );
  AOI222X1 U259 ( .IN1(data_csc[24]), .IN2(n653), .IN3(data_cot[24]), .IN4(
        n656), .IN5(data_sec[24]), .IN6(n660), .QN(n304) );
  AOI222X1 U260 ( .IN1(data_sin[24]), .IN2(n644), .IN3(data_tan[24]), .IN4(
        n650), .IN5(data_cos[24]), .IN6(n647), .QN(n303) );
  AOI222X1 U261 ( .IN1(data_csc[23]), .IN2(n652), .IN3(data_cot[23]), .IN4(
        n655), .IN5(data_sec[23]), .IN6(n659), .QN(n306) );
  AOI222X1 U262 ( .IN1(data_sin[23]), .IN2(n643), .IN3(data_tan[23]), .IN4(
        n650), .IN5(data_cos[23]), .IN6(n646), .QN(n305) );
  AOI222X1 U263 ( .IN1(data_csc[22]), .IN2(n652), .IN3(data_cot[22]), .IN4(
        n655), .IN5(data_sec[22]), .IN6(n659), .QN(n308) );
  AOI222X1 U264 ( .IN1(data_sin[22]), .IN2(n643), .IN3(data_tan[22]), .IN4(
        n650), .IN5(data_cos[22]), .IN6(n646), .QN(n307) );
  AOI222X1 U265 ( .IN1(data_csc[21]), .IN2(n652), .IN3(data_cot[21]), .IN4(
        n655), .IN5(data_sec[21]), .IN6(n659), .QN(n310) );
  AOI222X1 U266 ( .IN1(data_sin[21]), .IN2(n643), .IN3(data_tan[21]), .IN4(
        n650), .IN5(data_cos[21]), .IN6(n646), .QN(n309) );
  AOI222X1 U267 ( .IN1(data_csc[20]), .IN2(n652), .IN3(data_cot[20]), .IN4(
        n655), .IN5(data_sec[20]), .IN6(n659), .QN(n312) );
  AOI222X1 U268 ( .IN1(data_sin[20]), .IN2(n643), .IN3(data_tan[20]), .IN4(
        n650), .IN5(data_cos[20]), .IN6(n646), .QN(n311) );
  AOI222X1 U269 ( .IN1(data_csc[19]), .IN2(n652), .IN3(data_cot[19]), .IN4(
        n655), .IN5(data_sec[19]), .IN6(n659), .QN(n314) );
  AOI222X1 U270 ( .IN1(data_sin[19]), .IN2(n643), .IN3(data_tan[19]), .IN4(
        n650), .IN5(data_cos[19]), .IN6(n646), .QN(n313) );
  AOI222X1 U271 ( .IN1(data_csc[18]), .IN2(n652), .IN3(data_cot[18]), .IN4(
        n655), .IN5(data_sec[18]), .IN6(n659), .QN(n316) );
  AOI222X1 U272 ( .IN1(data_sin[18]), .IN2(n643), .IN3(data_tan[18]), .IN4(
        n650), .IN5(data_cos[18]), .IN6(n646), .QN(n315) );
  AOI222X1 U273 ( .IN1(data_csc[17]), .IN2(n652), .IN3(data_cot[17]), .IN4(
        n655), .IN5(data_sec[17]), .IN6(n659), .QN(n318) );
  AOI222X1 U274 ( .IN1(data_sin[17]), .IN2(n643), .IN3(data_tan[17]), .IN4(
        n650), .IN5(data_cos[17]), .IN6(n646), .QN(n317) );
  AOI222X1 U275 ( .IN1(data_csc[16]), .IN2(n652), .IN3(data_cot[16]), .IN4(
        n655), .IN5(data_sec[16]), .IN6(n659), .QN(n320) );
  AOI222X1 U276 ( .IN1(data_sin[16]), .IN2(n643), .IN3(data_tan[16]), .IN4(
        n650), .IN5(data_cos[16]), .IN6(n646), .QN(n319) );
  AOI222X1 U277 ( .IN1(data_csc[15]), .IN2(n652), .IN3(data_cot[15]), .IN4(
        n655), .IN5(data_sec[15]), .IN6(n659), .QN(n322) );
  AOI222X1 U278 ( .IN1(data_sin[15]), .IN2(n643), .IN3(data_tan[15]), .IN4(
        n650), .IN5(data_cos[15]), .IN6(n646), .QN(n321) );
  AOI222X1 U279 ( .IN1(data_csc[14]), .IN2(n652), .IN3(data_cot[14]), .IN4(
        n655), .IN5(data_sec[14]), .IN6(n659), .QN(n324) );
  AOI222X1 U280 ( .IN1(data_sin[14]), .IN2(n643), .IN3(data_tan[14]), .IN4(
        n650), .IN5(data_cos[14]), .IN6(n646), .QN(n323) );
  AOI222X1 U281 ( .IN1(data_csc[13]), .IN2(n652), .IN3(data_cot[13]), .IN4(
        n655), .IN5(data_sec[13]), .IN6(n659), .QN(n326) );
  AOI222X1 U282 ( .IN1(data_sin[13]), .IN2(n643), .IN3(data_tan[13]), .IN4(
        n650), .IN5(data_cos[13]), .IN6(n646), .QN(n325) );
  AOI222X1 U283 ( .IN1(data_csc[12]), .IN2(n652), .IN3(data_cot[12]), .IN4(
        n655), .IN5(data_sec[12]), .IN6(n659), .QN(n328) );
  AOI222X1 U284 ( .IN1(data_sin[12]), .IN2(n643), .IN3(data_tan[12]), .IN4(
        n650), .IN5(data_cos[12]), .IN6(n646), .QN(n327) );
  AOI222X1 U285 ( .IN1(data_csc[11]), .IN2(n651), .IN3(data_cot[11]), .IN4(
        n654), .IN5(data_sec[11]), .IN6(n658), .QN(n330) );
  AOI222X1 U286 ( .IN1(data_sin[11]), .IN2(n642), .IN3(data_tan[11]), .IN4(
        n650), .IN5(data_cos[11]), .IN6(n645), .QN(n329) );
  AOI222X1 U287 ( .IN1(data_csc[10]), .IN2(n651), .IN3(data_cot[10]), .IN4(
        n654), .IN5(data_sec[10]), .IN6(n658), .QN(n332) );
  AOI222X1 U288 ( .IN1(data_sin[10]), .IN2(n642), .IN3(data_tan[10]), .IN4(
        n650), .IN5(data_cos[10]), .IN6(n645), .QN(n331) );
  AOI222X1 U289 ( .IN1(data_csc[9]), .IN2(n651), .IN3(data_cot[9]), .IN4(n654), 
        .IN5(data_sec[9]), .IN6(n658), .QN(n334) );
  AOI222X1 U290 ( .IN1(data_sin[9]), .IN2(n642), .IN3(data_tan[9]), .IN4(n650), 
        .IN5(data_cos[9]), .IN6(n645), .QN(n333) );
  AOI222X1 U291 ( .IN1(data_csc[8]), .IN2(n651), .IN3(data_cot[8]), .IN4(n654), 
        .IN5(data_sec[8]), .IN6(n658), .QN(n336) );
  AOI222X1 U292 ( .IN1(data_sin[8]), .IN2(n642), .IN3(data_tan[8]), .IN4(n650), 
        .IN5(data_cos[8]), .IN6(n645), .QN(n335) );
  AOI222X1 U293 ( .IN1(data_csc[7]), .IN2(n651), .IN3(data_cot[7]), .IN4(n654), 
        .IN5(data_sec[7]), .IN6(n658), .QN(n338) );
  AOI222X1 U294 ( .IN1(data_sin[7]), .IN2(n642), .IN3(data_tan[7]), .IN4(n650), 
        .IN5(data_cos[7]), .IN6(n645), .QN(n337) );
  AOI222X1 U295 ( .IN1(data_csc[6]), .IN2(n651), .IN3(data_cot[6]), .IN4(n654), 
        .IN5(data_sec[6]), .IN6(n658), .QN(n340) );
  AOI222X1 U296 ( .IN1(data_sin[6]), .IN2(n642), .IN3(data_tan[6]), .IN4(n650), 
        .IN5(data_cos[6]), .IN6(n645), .QN(n339) );
  AOI222X1 U297 ( .IN1(data_csc[5]), .IN2(n651), .IN3(data_cot[5]), .IN4(n654), 
        .IN5(data_sec[5]), .IN6(n658), .QN(n342) );
  AOI222X1 U298 ( .IN1(data_sin[5]), .IN2(n642), .IN3(data_tan[5]), .IN4(n650), 
        .IN5(data_cos[5]), .IN6(n645), .QN(n341) );
  AOI222X1 U299 ( .IN1(data_csc[4]), .IN2(n651), .IN3(data_cot[4]), .IN4(n654), 
        .IN5(data_sec[4]), .IN6(n658), .QN(n344) );
  AOI222X1 U300 ( .IN1(data_sin[4]), .IN2(n642), .IN3(data_tan[4]), .IN4(n650), 
        .IN5(data_cos[4]), .IN6(n645), .QN(n343) );
  AOI222X1 U301 ( .IN1(data_csc[3]), .IN2(n651), .IN3(data_cot[3]), .IN4(n654), 
        .IN5(data_sec[3]), .IN6(n658), .QN(n346) );
  AOI222X1 U302 ( .IN1(data_sin[3]), .IN2(n642), .IN3(data_tan[3]), .IN4(n650), 
        .IN5(data_cos[3]), .IN6(n645), .QN(n345) );
  AOI222X1 U303 ( .IN1(data_csc[2]), .IN2(n651), .IN3(data_cot[2]), .IN4(n654), 
        .IN5(data_sec[2]), .IN6(n658), .QN(n348) );
  AOI222X1 U304 ( .IN1(data_sin[2]), .IN2(n642), .IN3(data_tan[2]), .IN4(n650), 
        .IN5(data_cos[2]), .IN6(n645), .QN(n347) );
  AOI222X1 U305 ( .IN1(data_csc[1]), .IN2(n651), .IN3(data_cot[1]), .IN4(n654), 
        .IN5(data_sec[1]), .IN6(n658), .QN(n350) );
  AOI222X1 U306 ( .IN1(data_sin[1]), .IN2(n642), .IN3(data_tan[1]), .IN4(n650), 
        .IN5(data_cos[1]), .IN6(n645), .QN(n349) );
  AOI222X1 U307 ( .IN1(data_csc[0]), .IN2(n651), .IN3(data_cot[0]), .IN4(n654), 
        .IN5(data_sec[0]), .IN6(n658), .QN(n352) );
  AOI222X1 U308 ( .IN1(data_sin[0]), .IN2(n642), .IN3(data_tan[0]), .IN4(n650), 
        .IN5(data_cos[0]), .IN6(n645), .QN(n351) );
  NAND3X0 U309 ( .IN1(actv[0]), .IN2(n823), .IN3(actv[2]), .QN(n354) );
  NAND3X0 U310 ( .IN1(n824), .IN2(n823), .IN3(actv[2]), .QN(n353) );
  NAND3X0 U311 ( .IN1(actv[0]), .IN2(n822), .IN3(actv[1]), .QN(n355) );
  OR3X1 U312 ( .IN1(n676), .IN2(n224), .IN3(n674), .Q(N357) );
  OR4X1 U313 ( .IN1(n672), .IN2(n676), .IN3(n670), .IN4(n668), .Q(N356) );
  AO22X1 U316 ( .IN1(N323), .IN2(n668), .IN3(degrees[31]), .IN4(n665), .Q(n368) );
  AO22X1 U318 ( .IN1(N91), .IN2(n676), .IN3(N124), .IN4(n674), .Q(n371) );
  OR2X1 U319 ( .IN1(n372), .IN2(n373), .Q(N354) );
  AO221X1 U320 ( .IN1(n666), .IN2(degrees_tmp1[30]), .IN3(N257), .IN4(n670), 
        .IN5(n374), .Q(n373) );
  AO22X1 U321 ( .IN1(N322), .IN2(n668), .IN3(degrees[30]), .IN4(n665), .Q(n374) );
  AO221X1 U322 ( .IN1(divider_out[30]), .IN2(n663), .IN3(N156), .IN4(n673), 
        .IN5(n375), .Q(n372) );
  AO22X1 U323 ( .IN1(N90), .IN2(n677), .IN3(N123), .IN4(n675), .Q(n375) );
  OR2X1 U324 ( .IN1(n376), .IN2(n377), .Q(N353) );
  AO221X1 U325 ( .IN1(n666), .IN2(degrees_tmp1[29]), .IN3(N256), .IN4(n670), 
        .IN5(n378), .Q(n377) );
  AO22X1 U326 ( .IN1(N321), .IN2(n668), .IN3(degrees[29]), .IN4(n665), .Q(n378) );
  AO221X1 U327 ( .IN1(divider_out[29]), .IN2(n663), .IN3(N155), .IN4(n673), 
        .IN5(n379), .Q(n376) );
  AO22X1 U328 ( .IN1(N89), .IN2(n677), .IN3(N122), .IN4(n675), .Q(n379) );
  OR2X1 U329 ( .IN1(n380), .IN2(n381), .Q(N352) );
  AO221X1 U330 ( .IN1(n666), .IN2(degrees_tmp1[28]), .IN3(N255), .IN4(n670), 
        .IN5(n382), .Q(n381) );
  AO22X1 U331 ( .IN1(N320), .IN2(n668), .IN3(degrees[28]), .IN4(n665), .Q(n382) );
  AO221X1 U332 ( .IN1(divider_out[28]), .IN2(n663), .IN3(N154), .IN4(n673), 
        .IN5(n383), .Q(n380) );
  AO22X1 U333 ( .IN1(N88), .IN2(n677), .IN3(N121), .IN4(n675), .Q(n383) );
  OR2X1 U334 ( .IN1(n384), .IN2(n385), .Q(N351) );
  AO221X1 U335 ( .IN1(n666), .IN2(degrees_tmp1[27]), .IN3(N254), .IN4(n670), 
        .IN5(n386), .Q(n385) );
  AO22X1 U336 ( .IN1(N319), .IN2(n668), .IN3(degrees[27]), .IN4(n665), .Q(n386) );
  AO221X1 U337 ( .IN1(divider_out[27]), .IN2(n663), .IN3(N153), .IN4(n673), 
        .IN5(n387), .Q(n384) );
  AO22X1 U338 ( .IN1(N87), .IN2(n677), .IN3(N120), .IN4(n675), .Q(n387) );
  OR2X1 U339 ( .IN1(n388), .IN2(n389), .Q(N350) );
  AO221X1 U340 ( .IN1(n666), .IN2(degrees_tmp1[26]), .IN3(N253), .IN4(n670), 
        .IN5(n390), .Q(n389) );
  AO22X1 U341 ( .IN1(N318), .IN2(n668), .IN3(degrees[26]), .IN4(n665), .Q(n390) );
  AO221X1 U342 ( .IN1(divider_out[26]), .IN2(n663), .IN3(N152), .IN4(n673), 
        .IN5(n391), .Q(n388) );
  AO22X1 U343 ( .IN1(N86), .IN2(n677), .IN3(N119), .IN4(n675), .Q(n391) );
  NAND3X0 U344 ( .IN1(n824), .IN2(n822), .IN3(actv[1]), .QN(n357) );
  OR2X1 U345 ( .IN1(n392), .IN2(n393), .Q(N349) );
  AO221X1 U346 ( .IN1(n666), .IN2(degrees_tmp1[25]), .IN3(N252), .IN4(n670), 
        .IN5(n394), .Q(n393) );
  AO22X1 U347 ( .IN1(N317), .IN2(n668), .IN3(degrees[25]), .IN4(n665), .Q(n394) );
  AO221X1 U348 ( .IN1(divider_out[25]), .IN2(n663), .IN3(N151), .IN4(n673), 
        .IN5(n395), .Q(n392) );
  AO22X1 U349 ( .IN1(N85), .IN2(n677), .IN3(N118), .IN4(n675), .Q(n395) );
  OR2X1 U350 ( .IN1(n396), .IN2(n397), .Q(N348) );
  AO221X1 U351 ( .IN1(n666), .IN2(degrees_tmp1[24]), .IN3(N251), .IN4(n670), 
        .IN5(n398), .Q(n397) );
  AO22X1 U352 ( .IN1(N316), .IN2(n668), .IN3(degrees[24]), .IN4(n665), .Q(n398) );
  AO221X1 U353 ( .IN1(divider_out[24]), .IN2(n663), .IN3(N150), .IN4(n672), 
        .IN5(n399), .Q(n396) );
  AO22X1 U354 ( .IN1(N84), .IN2(n677), .IN3(N117), .IN4(n674), .Q(n399) );
  OR2X1 U355 ( .IN1(n400), .IN2(n401), .Q(N347) );
  AO221X1 U356 ( .IN1(n666), .IN2(degrees_tmp1[23]), .IN3(N250), .IN4(n670), 
        .IN5(n402), .Q(n401) );
  AO22X1 U357 ( .IN1(N315), .IN2(n668), .IN3(degrees[23]), .IN4(n665), .Q(n402) );
  AO221X1 U358 ( .IN1(divider_out[23]), .IN2(n663), .IN3(N149), .IN4(n673), 
        .IN5(n403), .Q(n400) );
  AO22X1 U359 ( .IN1(N83), .IN2(n677), .IN3(N116), .IN4(n674), .Q(n403) );
  OR2X1 U360 ( .IN1(n404), .IN2(n405), .Q(N346) );
  AO221X1 U361 ( .IN1(n666), .IN2(degrees_tmp1[22]), .IN3(N249), .IN4(n670), 
        .IN5(n406), .Q(n405) );
  AO22X1 U362 ( .IN1(N314), .IN2(n668), .IN3(degrees[22]), .IN4(n665), .Q(n406) );
  AO221X1 U363 ( .IN1(divider_out[22]), .IN2(n663), .IN3(N148), .IN4(n673), 
        .IN5(n407), .Q(n404) );
  AO22X1 U364 ( .IN1(N82), .IN2(n677), .IN3(N115), .IN4(n674), .Q(n407) );
  OR2X1 U365 ( .IN1(n408), .IN2(n409), .Q(N345) );
  AO221X1 U366 ( .IN1(n666), .IN2(degrees_tmp1[21]), .IN3(N248), .IN4(n670), 
        .IN5(n410), .Q(n409) );
  AO22X1 U367 ( .IN1(N313), .IN2(n668), .IN3(degrees[21]), .IN4(n665), .Q(n410) );
  AO221X1 U368 ( .IN1(divider_out[21]), .IN2(n663), .IN3(N147), .IN4(n673), 
        .IN5(n411), .Q(n408) );
  AO22X1 U369 ( .IN1(N81), .IN2(n677), .IN3(N114), .IN4(n674), .Q(n411) );
  OR2X1 U370 ( .IN1(n412), .IN2(n413), .Q(N344) );
  AO221X1 U371 ( .IN1(n666), .IN2(degrees_tmp1[20]), .IN3(N247), .IN4(n670), 
        .IN5(n414), .Q(n413) );
  AO22X1 U372 ( .IN1(N312), .IN2(n668), .IN3(degrees[20]), .IN4(n665), .Q(n414) );
  AO221X1 U373 ( .IN1(divider_out[20]), .IN2(n663), .IN3(N146), .IN4(n672), 
        .IN5(n415), .Q(n412) );
  AO22X1 U374 ( .IN1(N80), .IN2(n677), .IN3(N113), .IN4(n674), .Q(n415) );
  OR2X1 U375 ( .IN1(n416), .IN2(n417), .Q(N343) );
  AO221X1 U376 ( .IN1(n667), .IN2(degrees_tmp1[19]), .IN3(N246), .IN4(n670), 
        .IN5(n418), .Q(n417) );
  AO22X1 U377 ( .IN1(N311), .IN2(n668), .IN3(degrees[19]), .IN4(n665), .Q(n418) );
  AO221X1 U378 ( .IN1(divider_out[19]), .IN2(n663), .IN3(N145), .IN4(n672), 
        .IN5(n419), .Q(n416) );
  AO22X1 U379 ( .IN1(N79), .IN2(n677), .IN3(N112), .IN4(n674), .Q(n419) );
  OR2X1 U380 ( .IN1(n420), .IN2(n421), .Q(N342) );
  AO221X1 U381 ( .IN1(n667), .IN2(degrees_tmp1[18]), .IN3(N245), .IN4(n670), 
        .IN5(n422), .Q(n421) );
  AO22X1 U382 ( .IN1(N310), .IN2(n668), .IN3(degrees[18]), .IN4(n664), .Q(n422) );
  AO221X1 U383 ( .IN1(divider_out[18]), .IN2(n663), .IN3(N144), .IN4(n672), 
        .IN5(n423), .Q(n420) );
  AO22X1 U384 ( .IN1(N78), .IN2(n677), .IN3(N111), .IN4(n674), .Q(n423) );
  OR2X1 U385 ( .IN1(n424), .IN2(n425), .Q(N341) );
  AO221X1 U386 ( .IN1(n667), .IN2(degrees_tmp1[17]), .IN3(N244), .IN4(n670), 
        .IN5(n426), .Q(n425) );
  AO22X1 U387 ( .IN1(N309), .IN2(n668), .IN3(degrees[17]), .IN4(n664), .Q(n426) );
  AO221X1 U388 ( .IN1(divider_out[17]), .IN2(n663), .IN3(N143), .IN4(n672), 
        .IN5(n427), .Q(n424) );
  AO22X1 U389 ( .IN1(N77), .IN2(n677), .IN3(N110), .IN4(n674), .Q(n427) );
  OR2X1 U390 ( .IN1(n428), .IN2(n429), .Q(N340) );
  AO221X1 U391 ( .IN1(n667), .IN2(degrees_tmp1[16]), .IN3(N243), .IN4(n670), 
        .IN5(n430), .Q(n429) );
  AO22X1 U392 ( .IN1(N308), .IN2(n668), .IN3(degrees[16]), .IN4(n664), .Q(n430) );
  AO221X1 U393 ( .IN1(divider_out[16]), .IN2(n663), .IN3(N142), .IN4(n672), 
        .IN5(n431), .Q(n428) );
  AO22X1 U394 ( .IN1(N76), .IN2(n677), .IN3(N109), .IN4(n674), .Q(n431) );
  NAND3X0 U395 ( .IN1(n823), .IN2(n822), .IN3(actv[0]), .QN(n356) );
  OR2X1 U396 ( .IN1(n432), .IN2(n433), .Q(N339) );
  AO221X1 U397 ( .IN1(n667), .IN2(degrees_tmp1[15]), .IN3(N242), .IN4(n671), 
        .IN5(n434), .Q(n433) );
  AO22X1 U398 ( .IN1(N307), .IN2(n668), .IN3(degrees[15]), .IN4(n664), .Q(n434) );
  AO221X1 U399 ( .IN1(divider_out[15]), .IN2(n663), .IN3(N141), .IN4(n672), 
        .IN5(n435), .Q(n432) );
  AO22X1 U400 ( .IN1(N75), .IN2(n676), .IN3(N108), .IN4(n674), .Q(n435) );
  OR2X1 U401 ( .IN1(n436), .IN2(n437), .Q(N338) );
  AO221X1 U402 ( .IN1(n667), .IN2(degrees_tmp1[14]), .IN3(N241), .IN4(n671), 
        .IN5(n438), .Q(n437) );
  AO22X1 U403 ( .IN1(N306), .IN2(n668), .IN3(degrees[14]), .IN4(n664), .Q(n438) );
  AO221X1 U404 ( .IN1(divider_out[14]), .IN2(n663), .IN3(N140), .IN4(n672), 
        .IN5(n439), .Q(n436) );
  AO22X1 U405 ( .IN1(N74), .IN2(n676), .IN3(N107), .IN4(n674), .Q(n439) );
  OR2X1 U406 ( .IN1(n440), .IN2(n441), .Q(N337) );
  AO221X1 U407 ( .IN1(n667), .IN2(degrees_tmp1[13]), .IN3(N240), .IN4(n671), 
        .IN5(n442), .Q(n441) );
  AO22X1 U408 ( .IN1(N305), .IN2(n668), .IN3(degrees[13]), .IN4(n664), .Q(n442) );
  AO221X1 U409 ( .IN1(divider_out[13]), .IN2(n663), .IN3(N139), .IN4(n672), 
        .IN5(n443), .Q(n440) );
  AO22X1 U410 ( .IN1(N73), .IN2(n676), .IN3(N106), .IN4(n674), .Q(n443) );
  OR2X1 U411 ( .IN1(n444), .IN2(n445), .Q(N336) );
  AO221X1 U412 ( .IN1(n667), .IN2(degrees_tmp1[12]), .IN3(N239), .IN4(n671), 
        .IN5(n446), .Q(n445) );
  AO22X1 U413 ( .IN1(N304), .IN2(n668), .IN3(degrees[12]), .IN4(n664), .Q(n446) );
  AO221X1 U414 ( .IN1(divider_out[12]), .IN2(n662), .IN3(N138), .IN4(n672), 
        .IN5(n447), .Q(n444) );
  AO22X1 U415 ( .IN1(N72), .IN2(n676), .IN3(N105), .IN4(n674), .Q(n447) );
  OR2X1 U416 ( .IN1(n448), .IN2(n449), .Q(N335) );
  AO221X1 U417 ( .IN1(n667), .IN2(degrees_tmp1[11]), .IN3(N238), .IN4(n671), 
        .IN5(n450), .Q(n449) );
  AO22X1 U418 ( .IN1(N303), .IN2(n669), .IN3(degrees[11]), .IN4(n664), .Q(n450) );
  AO221X1 U419 ( .IN1(divider_out[11]), .IN2(n662), .IN3(N137), .IN4(n672), 
        .IN5(n451), .Q(n448) );
  AO22X1 U420 ( .IN1(N71), .IN2(n676), .IN3(N104), .IN4(n674), .Q(n451) );
  OR2X1 U421 ( .IN1(n452), .IN2(n453), .Q(N334) );
  AO221X1 U422 ( .IN1(n667), .IN2(degrees_tmp1[10]), .IN3(N237), .IN4(n671), 
        .IN5(n454), .Q(n453) );
  AO22X1 U423 ( .IN1(N302), .IN2(n669), .IN3(degrees[10]), .IN4(n664), .Q(n454) );
  AO221X1 U424 ( .IN1(divider_out[10]), .IN2(n662), .IN3(N136), .IN4(n672), 
        .IN5(n455), .Q(n452) );
  AO22X1 U425 ( .IN1(N70), .IN2(n676), .IN3(N103), .IN4(n674), .Q(n455) );
  OR2X1 U426 ( .IN1(n456), .IN2(n457), .Q(N333) );
  AO221X1 U427 ( .IN1(n667), .IN2(degrees_tmp1[9]), .IN3(N236), .IN4(n671), 
        .IN5(n458), .Q(n457) );
  AO22X1 U428 ( .IN1(N301), .IN2(n669), .IN3(degrees[9]), .IN4(n664), .Q(n458)
         );
  AO221X1 U429 ( .IN1(divider_out[9]), .IN2(n662), .IN3(N135), .IN4(n672), 
        .IN5(n459), .Q(n456) );
  AO22X1 U430 ( .IN1(N69), .IN2(n676), .IN3(N102), .IN4(n674), .Q(n459) );
  OR2X1 U431 ( .IN1(n460), .IN2(n461), .Q(N332) );
  AO221X1 U432 ( .IN1(n667), .IN2(degrees_tmp1[8]), .IN3(N235), .IN4(n671), 
        .IN5(n462), .Q(n461) );
  AO22X1 U433 ( .IN1(N300), .IN2(n669), .IN3(n664), .IN4(degrees[8]), .Q(n462)
         );
  AO221X1 U434 ( .IN1(N101), .IN2(n675), .IN3(N68), .IN4(n676), .IN5(n463), 
        .Q(n460) );
  AO22X1 U435 ( .IN1(N134), .IN2(n673), .IN3(n662), .IN4(divider_out[8]), .Q(
        n463) );
  OR2X1 U436 ( .IN1(n464), .IN2(n465), .Q(N331) );
  AO221X1 U437 ( .IN1(n667), .IN2(degrees_tmp1[7]), .IN3(N234), .IN4(n671), 
        .IN5(n466), .Q(n465) );
  AO22X1 U438 ( .IN1(N299), .IN2(n669), .IN3(n665), .IN4(degrees[7]), .Q(n466)
         );
  AO221X1 U439 ( .IN1(N100), .IN2(n675), .IN3(N67), .IN4(n676), .IN5(n467), 
        .Q(n464) );
  AO22X1 U440 ( .IN1(N133), .IN2(n673), .IN3(n662), .IN4(divider_out[7]), .Q(
        n467) );
  OR2X1 U441 ( .IN1(n468), .IN2(n469), .Q(N330) );
  AO221X1 U442 ( .IN1(n666), .IN2(degrees_tmp1[6]), .IN3(N233), .IN4(n671), 
        .IN5(n470), .Q(n469) );
  AO22X1 U443 ( .IN1(N298), .IN2(n669), .IN3(n664), .IN4(degrees[6]), .Q(n470)
         );
  AO221X1 U444 ( .IN1(divider_out[6]), .IN2(n662), .IN3(N132), .IN4(n672), 
        .IN5(n471), .Q(n468) );
  AO22X1 U445 ( .IN1(N66), .IN2(n676), .IN3(N99), .IN4(n674), .Q(n471) );
  NAND3X0 U446 ( .IN1(n823), .IN2(n822), .IN3(n824), .QN(n358) );
  OR2X1 U447 ( .IN1(n472), .IN2(n473), .Q(N329) );
  AO221X1 U448 ( .IN1(n667), .IN2(degrees_tmp1[5]), .IN3(N232), .IN4(n671), 
        .IN5(n474), .Q(n473) );
  AO22X1 U449 ( .IN1(N297), .IN2(n669), .IN3(n665), .IN4(degrees[5]), .Q(n474)
         );
  AO221X1 U450 ( .IN1(N98), .IN2(n675), .IN3(N65), .IN4(n676), .IN5(n475), .Q(
        n472) );
  AO22X1 U451 ( .IN1(N131), .IN2(n673), .IN3(n662), .IN4(divider_out[5]), .Q(
        n475) );
  OR2X1 U452 ( .IN1(n476), .IN2(n477), .Q(N328) );
  AO221X1 U453 ( .IN1(n666), .IN2(degrees_tmp1[4]), .IN3(N231), .IN4(n671), 
        .IN5(n478), .Q(n477) );
  AO22X1 U454 ( .IN1(N296), .IN2(n669), .IN3(n664), .IN4(degrees[4]), .Q(n478)
         );
  AO221X1 U455 ( .IN1(N97), .IN2(n675), .IN3(N64), .IN4(n676), .IN5(n479), .Q(
        n476) );
  AO22X1 U456 ( .IN1(N130), .IN2(n673), .IN3(n662), .IN4(divider_out[4]), .Q(
        n479) );
  OR2X1 U457 ( .IN1(n480), .IN2(n481), .Q(N327) );
  AO221X1 U458 ( .IN1(n667), .IN2(degrees_tmp1[3]), .IN3(N230), .IN4(n671), 
        .IN5(n482), .Q(n481) );
  AO22X1 U459 ( .IN1(N295), .IN2(n669), .IN3(n665), .IN4(degrees[3]), .Q(n482)
         );
  AO221X1 U460 ( .IN1(N96), .IN2(n675), .IN3(N63), .IN4(n676), .IN5(n483), .Q(
        n480) );
  AO22X1 U461 ( .IN1(N129), .IN2(n673), .IN3(n662), .IN4(divider_out[3]), .Q(
        n483) );
  OR2X1 U462 ( .IN1(n484), .IN2(n485), .Q(N326) );
  AO221X1 U463 ( .IN1(n666), .IN2(degrees_tmp1[2]), .IN3(N229), .IN4(n671), 
        .IN5(n486), .Q(n485) );
  AO22X1 U464 ( .IN1(N294), .IN2(n669), .IN3(n664), .IN4(degrees[2]), .Q(n486)
         );
  AO221X1 U465 ( .IN1(N95), .IN2(n675), .IN3(N62), .IN4(n676), .IN5(n487), .Q(
        n484) );
  OR2X1 U467 ( .IN1(n488), .IN2(n489), .Q(N325) );
  AO221X1 U468 ( .IN1(n667), .IN2(n639), .IN3(N228), .IN4(n671), .IN5(n490), 
        .Q(n489) );
  AO22X1 U469 ( .IN1(N293), .IN2(n669), .IN3(degrees[1]), .IN4(n664), .Q(n490)
         );
  AO221X1 U470 ( .IN1(N94), .IN2(n675), .IN3(N61), .IN4(n676), .IN5(n491), .Q(
        n488) );
  OR2X1 U472 ( .IN1(n492), .IN2(n493), .Q(N324) );
  AO221X1 U473 ( .IN1(n666), .IN2(degrees_tmp1[0]), .IN3(N227), .IN4(n671), 
        .IN5(n494), .Q(n493) );
  AO22X1 U474 ( .IN1(N292), .IN2(n669), .IN3(degrees[0]), .IN4(n664), .Q(n494)
         );
  AO21X1 U477 ( .IN1(n498), .IN2(n499), .IN3(N44), .Q(n497) );
  OR4X1 U478 ( .IN1(degrees[28]), .IN2(degrees[29]), .IN3(degrees[30]), .IN4(
        degrees[31]), .Q(n501) );
  OR4X1 U479 ( .IN1(degrees[3]), .IN2(degrees[6]), .IN3(degrees[8]), .IN4(
        degrees[9]), .Q(n500) );
  NAND4X0 U480 ( .IN1(degrees[7]), .IN2(degrees[4]), .IN3(degrees[2]), .IN4(
        degrees[5]), .QN(n507) );
  AO21X1 U482 ( .IN1(n509), .IN2(n510), .IN3(N41), .Q(n508) );
  NAND4X0 U483 ( .IN1(n806), .IN2(n805), .IN3(n804), .IN4(n803), .QN(n503) );
  NAND4X0 U484 ( .IN1(n802), .IN2(n801), .IN3(n800), .IN4(n799), .QN(n502) );
  OR4X1 U485 ( .IN1(degrees[28]), .IN2(degrees[29]), .IN3(degrees[2]), .IN4(
        degrees[30]), .Q(n512) );
  OR4X1 U486 ( .IN1(degrees[31]), .IN2(degrees[4]), .IN3(degrees[7]), .IN4(
        degrees[9]), .Q(n511) );
  NAND4X0 U487 ( .IN1(degrees[8]), .IN2(degrees[6]), .IN3(degrees[5]), .IN4(
        degrees[3]), .QN(n513) );
  NAND4X0 U488 ( .IN1(n818), .IN2(n816), .IN3(n815), .IN4(n814), .QN(n506) );
  NAND4X0 U489 ( .IN1(n813), .IN2(n812), .IN3(n811), .IN4(n810), .QN(n505) );
  NAND4X0 U490 ( .IN1(n809), .IN2(n808), .IN3(n807), .IN4(n817), .QN(n504) );
  AO221X1 U491 ( .IN1(divider_out[0]), .IN2(n662), .IN3(N126), .IN4(n673), 
        .IN5(n514), .Q(n492) );
  AO21X1 U495 ( .IN1(n518), .IN2(n519), .IN3(N52), .Q(n517) );
  OR4X1 U496 ( .IN1(divider_out[21]), .IN2(divider_out[22]), .IN3(
        divider_out[23]), .IN4(divider_out[24]), .Q(n523) );
  OR4X1 U497 ( .IN1(divider_out[25]), .IN2(divider_out[26]), .IN3(
        divider_out[27]), .IN4(divider_out[28]), .Q(n522) );
  OR4X1 U498 ( .IN1(divider_out[29]), .IN2(divider_out[30]), .IN3(
        divider_out[31]), .IN4(divider_out[4]), .Q(n521) );
  OR4X1 U499 ( .IN1(divider_out[5]), .IN2(divider_out[6]), .IN3(divider_out[7]), .IN4(divider_out[9]), .Q(n520) );
  OR4X1 U501 ( .IN1(divider_out[17]), .IN2(divider_out[18]), .IN3(
        divider_out[19]), .IN4(divider_out[20]), .Q(n524) );
  AO21X1 U502 ( .IN1(n529), .IN2(n530), .IN3(N55), .Q(n528) );
  OR4X1 U503 ( .IN1(divider_out[20]), .IN2(divider_out[21]), .IN3(
        divider_out[22]), .IN4(divider_out[23]), .Q(n534) );
  OR4X1 U504 ( .IN1(divider_out[24]), .IN2(divider_out[25]), .IN3(
        divider_out[26]), .IN4(divider_out[27]), .Q(n533) );
  OR4X1 U505 ( .IN1(divider_out[28]), .IN2(divider_out[29]), .IN3(
        divider_out[30]), .IN4(divider_out[31]), .Q(n532) );
  OR4X1 U506 ( .IN1(divider_out[3]), .IN2(divider_out[6]), .IN3(divider_out[8]), .IN4(divider_out[9]), .Q(n531) );
  NAND4X0 U507 ( .IN1(divider_out[7]), .IN2(divider_out[5]), .IN3(
        divider_out[4]), .IN4(divider_out[2]), .QN(n536) );
  NAND4X0 U508 ( .IN1(n796), .IN2(n795), .IN3(n794), .IN4(n793), .QN(n526) );
  NAND4X0 U509 ( .IN1(n792), .IN2(n791), .IN3(n790), .IN4(n789), .QN(n525) );
  sine_lut a1 ( .quad(quad), .enable(sin_enable), .degrees(degrees_tmp2), 
        .data({data_sin[63], SYNOPSYS_UNCONNECTED__0, data_sin[61:0]}), .rst(
        rst), .clk(clk) );
  cosine_lut a2 ( .quad(quad), .enable(cos_enable), .degrees(degrees_tmp2), 
        .data({data_cos[63], SYNOPSYS_UNCONNECTED__1, data_cos[61:0]}), .rst(
        rst), .clk(clk) );
  tangent_lut a3 ( .quad(quad), .enable(tan_enable), .degrees(degrees_tmp2), 
        .data(data_tan), .rst(rst), .clk(clk) );
  cosecant_lut a4 ( .quad(quad), .enable(csc_enable), .degrees(degrees_tmp2), 
        .data(data_csc), .rst(rst), .clk(clk) );
  secant_lut a5 ( .quad(quad), .enable(sec_enable), .degrees(degrees_tmp2), 
        .data(data_sec), .rst(rst), .clk(clk) );
  cotangent_lut a6 ( .quad(quad), .enable(cot_enable), .degrees(degrees_tmp2), 
        .data(data_cot), .rst(rst), .clk(clk) );
  dividor a7 ( .clk(clk), .inp(degrees), .rst(rst), .out(divider_out) );
  top_DW01_sub_0 sub_187 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0}), .B(degrees), .CI(1'b0), .DIFF({N323, N322, N321, N320, N319, N318, N317, 
        N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, 
        N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, 
        N292}) );
  top_DW01_sub_1 sub_168 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0}), .B({degrees_tmp1[31:2], n639, degrees_tmp1[0]}), .CI(1'b0), .DIFF({N258, 
        N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, 
        N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, 
        N233, N232, N231, N230, N229, N228, N227}) );
  top_DW01_sub_2 sub_162 ( .A(degrees), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 
        1'b0, 1'b0}), .CI(1'b0), .DIFF({N224, N223, N222, N221, N220, N219, 
        N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, 
        N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, 
        N194, N193}) );
  top_DW01_sub_3 sub_144 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0}), .B(divider_out), .CI(1'b0), .DIFF({N157, N156, N155, N154, N153, N152, N151, 
        N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, 
        N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, 
        N126}) );
  top_DW01_sub_4 sub_138 ( .A(divider_out), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 
        1'b1, 1'b0, 1'b0}), .CI(1'b0), .DIFF({N124, N123, N122, N121, N120, 
        N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, 
        N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, 
        N95, N94, N93}) );
  top_DW01_sub_5 sub_131 ( .A(divider_out), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        1'b1, 1'b1, 1'b0}), .CI(1'b0), .DIFF({N91, N90, N89, N88, N87, N86, 
        N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, 
        N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60}) );
  DFFX1 \degrees_tmp1_reg[6]  ( .D(n543), .CLK(clk), .Q(degrees_tmp1[6]) );
  DFFX1 \degrees_tmp1_reg[4]  ( .D(n541), .CLK(clk), .Q(degrees_tmp1[4]) );
  DFFX1 \degrees_tmp1_reg[2]  ( .D(n539), .CLK(clk), .Q(degrees_tmp1[2]) );
  DFFX1 \degrees_tmp1_reg[29]  ( .D(n566), .CLK(clk), .Q(degrees_tmp1[29]) );
  DFFX1 \degrees_tmp1_reg[23]  ( .D(n560), .CLK(clk), .Q(degrees_tmp1[23]) );
  DFFX1 \degrees_tmp1_reg[17]  ( .D(n554), .CLK(clk), .Q(degrees_tmp1[17]) );
  DFFX1 \degrees_tmp1_reg[11]  ( .D(n548), .CLK(clk), .Q(degrees_tmp1[11]) );
  DFFX1 \degrees_tmp1_reg[28]  ( .D(n565), .CLK(clk), .Q(degrees_tmp1[28]) );
  DFFX1 \degrees_tmp1_reg[22]  ( .D(n559), .CLK(clk), .Q(degrees_tmp1[22]) );
  DFFX1 \degrees_tmp1_reg[16]  ( .D(n553), .CLK(clk), .Q(degrees_tmp1[16]) );
  DFFX1 \degrees_tmp1_reg[10]  ( .D(n547), .CLK(clk), .Q(degrees_tmp1[10]) );
  DFFX1 \degrees_tmp1_reg[27]  ( .D(n564), .CLK(clk), .Q(degrees_tmp1[27]) );
  DFFX1 \degrees_tmp1_reg[21]  ( .D(n558), .CLK(clk), .Q(degrees_tmp1[21]) );
  DFFX1 \degrees_tmp1_reg[15]  ( .D(n552), .CLK(clk), .Q(degrees_tmp1[15]) );
  DFFX1 \degrees_tmp1_reg[30]  ( .D(n567), .CLK(clk), .Q(degrees_tmp1[30]) );
  DFFX1 \degrees_tmp1_reg[26]  ( .D(n563), .CLK(clk), .Q(degrees_tmp1[26]) );
  DFFX1 \degrees_tmp1_reg[20]  ( .D(n557), .CLK(clk), .Q(degrees_tmp1[20]) );
  DFFX1 \degrees_tmp1_reg[14]  ( .D(n551), .CLK(clk), .Q(degrees_tmp1[14]) );
  DFFX1 \degrees_tmp1_reg[24]  ( .D(n561), .CLK(clk), .Q(degrees_tmp1[24]) );
  DFFX1 \degrees_tmp1_reg[18]  ( .D(n555), .CLK(clk), .Q(degrees_tmp1[18]) );
  DFFX1 \degrees_tmp1_reg[12]  ( .D(n549), .CLK(clk), .Q(degrees_tmp1[12]) );
  DFFX1 \degrees_tmp1_reg[9]  ( .D(n546), .CLK(clk), .Q(degrees_tmp1[9]) );
  DFFX1 \degrees_tmp1_reg[8]  ( .D(n545), .CLK(clk), .Q(degrees_tmp1[8]) );
  DFFX1 \degrees_tmp1_reg[25]  ( .D(n562), .CLK(clk), .Q(degrees_tmp1[25]) );
  DFFX1 \degrees_tmp1_reg[19]  ( .D(n556), .CLK(clk), .Q(degrees_tmp1[19]) );
  DFFX1 \degrees_tmp1_reg[13]  ( .D(n550), .CLK(clk), .Q(degrees_tmp1[13]) );
  DFFX1 \degrees_tmp1_reg[7]  ( .D(n544), .CLK(clk), .Q(degrees_tmp1[7]), .QN(
        n694) );
  DFFX1 \degrees_tmp1_reg[5]  ( .D(n542), .CLK(clk), .Q(degrees_tmp1[5]), .QN(
        n693) );
  DFFX1 \degrees_tmp1_reg[31]  ( .D(n568), .CLK(clk), .Q(degrees_tmp1[31]) );
  DFFX1 \degrees_tmp1_reg[3]  ( .D(n540), .CLK(clk), .Q(degrees_tmp1[3]) );
  DFFX1 \degrees_tmp1_reg[0]  ( .D(n537), .CLK(clk), .Q(degrees_tmp1[0]) );
  DFFX1 \data1_reg[61]  ( .D(N445), .CLK(clk), .Q(data1[61]) );
  DFFX1 \data1_reg[60]  ( .D(N444), .CLK(clk), .Q(data1[60]) );
  DFFX1 \data1_reg[59]  ( .D(N443), .CLK(clk), .Q(data1[59]) );
  DFFX1 \data1_reg[58]  ( .D(N442), .CLK(clk), .Q(data1[58]) );
  DFFX1 \data1_reg[57]  ( .D(N441), .CLK(clk), .Q(data1[57]) );
  DFFX1 \data1_reg[56]  ( .D(N440), .CLK(clk), .Q(data1[56]) );
  DFFX1 \data1_reg[55]  ( .D(N439), .CLK(clk), .Q(data1[55]) );
  DFFX1 \data1_reg[54]  ( .D(N438), .CLK(clk), .Q(data1[54]) );
  DFFX1 \data1_reg[53]  ( .D(N437), .CLK(clk), .Q(data1[53]) );
  DFFX1 \data1_reg[50]  ( .D(N434), .CLK(clk), .Q(data1[50]) );
  DFFX1 \data1_reg[49]  ( .D(N433), .CLK(clk), .Q(data1[49]) );
  DFFX1 \data1_reg[48]  ( .D(N432), .CLK(clk), .Q(data1[48]) );
  DFFX1 \data1_reg[47]  ( .D(N431), .CLK(clk), .Q(data1[47]) );
  DFFX1 \data1_reg[46]  ( .D(N430), .CLK(clk), .Q(data1[46]) );
  DFFX1 \data1_reg[45]  ( .D(N429), .CLK(clk), .Q(data1[45]) );
  DFFX1 \data1_reg[44]  ( .D(N428), .CLK(clk), .Q(data1[44]) );
  DFFX1 \data1_reg[43]  ( .D(N427), .CLK(clk), .Q(data1[43]) );
  DFFX1 \data1_reg[42]  ( .D(N426), .CLK(clk), .Q(data1[42]) );
  DFFX1 \data1_reg[41]  ( .D(N425), .CLK(clk), .Q(data1[41]) );
  DFFX1 \data1_reg[40]  ( .D(N424), .CLK(clk), .Q(data1[40]) );
  DFFX1 \data1_reg[39]  ( .D(N423), .CLK(clk), .Q(data1[39]) );
  DFFX1 \data1_reg[38]  ( .D(N422), .CLK(clk), .Q(data1[38]) );
  DFFX1 \data1_reg[37]  ( .D(N421), .CLK(clk), .Q(data1[37]) );
  DFFX1 \data1_reg[36]  ( .D(N420), .CLK(clk), .Q(data1[36]) );
  DFFX1 \data1_reg[35]  ( .D(N419), .CLK(clk), .Q(data1[35]) );
  DFFX1 \data1_reg[34]  ( .D(N418), .CLK(clk), .Q(data1[34]) );
  DFFX1 \data1_reg[33]  ( .D(N417), .CLK(clk), .Q(data1[33]) );
  DFFX1 \data1_reg[32]  ( .D(N416), .CLK(clk), .Q(data1[32]) );
  DFFX1 \data1_reg[31]  ( .D(N415), .CLK(clk), .Q(data1[31]) );
  DFFX1 \data1_reg[30]  ( .D(N414), .CLK(clk), .Q(data1[30]) );
  DFFX1 \data1_reg[29]  ( .D(N413), .CLK(clk), .Q(data1[29]) );
  DFFX1 \data1_reg[28]  ( .D(N412), .CLK(clk), .Q(data1[28]) );
  DFFX1 \data1_reg[27]  ( .D(N411), .CLK(clk), .Q(data1[27]) );
  INVX0 U511 ( .INP(n496), .ZN(n798) );
  INVX0 U512 ( .INP(n631), .ZN(n676) );
  INVX0 U513 ( .INP(n631), .ZN(n677) );
  INVX0 U514 ( .INP(n224), .ZN(n679) );
  INVX0 U515 ( .INP(n633), .ZN(n668) );
  INVX0 U516 ( .INP(n632), .ZN(n665) );
  INVX0 U517 ( .INP(n632), .ZN(n664) );
  INVX0 U518 ( .INP(n633), .ZN(n669) );
  INVX0 U519 ( .INP(n358), .ZN(n642) );
  INVX0 U520 ( .INP(n358), .ZN(n643) );
  INVX0 U521 ( .INP(n358), .ZN(n644) );
  INVX0 U522 ( .INP(n634), .ZN(n674) );
  INVX0 U523 ( .INP(n636), .ZN(n673) );
  INVX0 U524 ( .INP(n634), .ZN(n675) );
  INVX0 U525 ( .INP(n635), .ZN(n662) );
  INVX0 U526 ( .INP(n516), .ZN(n788) );
  INVX0 U527 ( .INP(n638), .ZN(n670) );
  INVX0 U528 ( .INP(n636), .ZN(n672) );
  INVX0 U529 ( .INP(n638), .ZN(n671) );
  INVX0 U530 ( .INP(n637), .ZN(n667) );
  INVX0 U531 ( .INP(n637), .ZN(n666) );
  INVX0 U532 ( .INP(n635), .ZN(n663) );
  OR2X1 U533 ( .IN1(n787), .IN2(n797), .Q(n631) );
  INVX0 U534 ( .INP(n357), .ZN(n649) );
  INVX0 U535 ( .INP(n357), .ZN(n650) );
  INVX0 U536 ( .INP(n353), .ZN(n658) );
  INVX0 U537 ( .INP(n356), .ZN(n645) );
  INVX0 U538 ( .INP(n353), .ZN(n659) );
  INVX0 U539 ( .INP(n356), .ZN(n646) );
  INVX0 U540 ( .INP(n353), .ZN(n660) );
  INVX0 U541 ( .INP(n356), .ZN(n647) );
  INVX0 U542 ( .INP(n353), .ZN(n661) );
  INVX0 U543 ( .INP(n356), .ZN(n648) );
  INVX0 U544 ( .INP(n354), .ZN(n654) );
  INVX0 U545 ( .INP(n354), .ZN(n655) );
  INVX0 U546 ( .INP(n354), .ZN(n656) );
  INVX0 U547 ( .INP(n354), .ZN(n657) );
  INVX0 U548 ( .INP(n355), .ZN(n651) );
  INVX0 U549 ( .INP(n355), .ZN(n652) );
  INVX0 U550 ( .INP(n355), .ZN(n653) );
  NAND3X0 U551 ( .IN1(n495), .IN2(n797), .IN3(n496), .QN(n632) );
  NAND3X0 U552 ( .IN1(n495), .IN2(n797), .IN3(n798), .QN(n633) );
  INVX0 U553 ( .INP(n358), .ZN(n820) );
  NBUFFX2 U554 ( .INP(n224), .Z(n678) );
  INVX0 U555 ( .INP(n732), .ZN(n741) );
  INVX0 U556 ( .INP(n735), .ZN(n740) );
  NAND2X1 U557 ( .IN1(N51), .IN2(n517), .QN(n516) );
  NOR4X0 U558 ( .IN1(n524), .IN2(n525), .IN3(n526), .IN4(n527), .QN(n518) );
  NAND3X0 U559 ( .IN1(N39), .IN2(n787), .IN3(n788), .QN(n634) );
  AO22X1 U560 ( .IN1(N127), .IN2(n673), .IN3(n662), .IN4(divider_out[1]), .Q(
        n491) );
  NAND4X0 U561 ( .IN1(N39), .IN2(n515), .IN3(n516), .IN4(n787), .QN(n635) );
  OR4X1 U562 ( .IN1(n515), .IN2(n797), .IN3(n788), .IN4(N50), .Q(n636) );
  OR2X1 U563 ( .IN1(n679), .IN2(N225), .Q(n637) );
  INVX0 U564 ( .INP(N50), .ZN(n787) );
  NAND2X1 U565 ( .IN1(N225), .IN2(n224), .QN(n638) );
  INVX0 U566 ( .INP(N39), .ZN(n797) );
  NAND2X1 U567 ( .IN1(N40), .IN2(n508), .QN(n495) );
  NOR4X0 U568 ( .IN1(n511), .IN2(n512), .IN3(n502), .IN4(n503), .QN(n510) );
  NOR2X0 U569 ( .IN1(n495), .IN2(N39), .QN(n224) );
  NOR2X0 U570 ( .IN1(n356), .IN2(n359), .QN(N34) );
  NOR2X0 U571 ( .IN1(n358), .IN2(n359), .QN(N33) );
  NOR2X0 U572 ( .IN1(n354), .IN2(n359), .QN(N38) );
  NOR2X0 U573 ( .IN1(n355), .IN2(n359), .QN(N36) );
  NOR2X0 U574 ( .IN1(n353), .IN2(n359), .QN(N37) );
  NOR2X0 U575 ( .IN1(n357), .IN2(n359), .QN(N35) );
  NAND2X1 U576 ( .IN1(N43), .IN2(n497), .QN(n496) );
  NOR4X0 U577 ( .IN1(n500), .IN2(n501), .IN3(n502), .IN4(n503), .QN(n499) );
  INVX0 U578 ( .INP(n355), .ZN(n821) );
  AND3X1 U579 ( .IN1(divider_out[2]), .IN2(divider_out[1]), .IN3(
        divider_out[3]), .Q(n752) );
  INVX0 U580 ( .INP(divider_out[7]), .ZN(n708) );
  NAND3X0 U581 ( .IN1(divider_out[1]), .IN2(divider_out[0]), .IN3(
        divider_out[3]), .QN(n695) );
  AO22X1 U582 ( .IN1(N60), .IN2(n677), .IN3(N93), .IN4(n675), .Q(n514) );
  AO22X1 U583 ( .IN1(N128), .IN2(n673), .IN3(n662), .IN4(divider_out[2]), .Q(
        n487) );
  NAND2X1 U584 ( .IN1(N54), .IN2(n528), .QN(n515) );
  INVX0 U585 ( .INP(divider_out[10]), .ZN(n795) );
  INVX0 U586 ( .INP(divider_out[11]), .ZN(n794) );
  INVX0 U587 ( .INP(divider_out[13]), .ZN(n792) );
  INVX0 U588 ( .INP(divider_out[14]), .ZN(n791) );
  INVX0 U589 ( .INP(divider_out[15]), .ZN(n790) );
  NAND3X0 U590 ( .IN1(n639), .IN2(degrees_tmp1[0]), .IN3(degrees_tmp1[3]), 
        .QN(n680) );
  INVX0 U591 ( .INP(divider_out[5]), .ZN(n739) );
  INVX0 U592 ( .INP(divider_out[4]), .ZN(n738) );
  INVX0 U593 ( .INP(divider_out[12]), .ZN(n793) );
  INVX0 U594 ( .INP(divider_out[16]), .ZN(n789) );
  NOR4X0 U595 ( .IN1(n535), .IN2(n525), .IN3(n526), .IN4(n536), .QN(n529) );
  OR4X1 U596 ( .IN1(divider_out[17]), .IN2(divider_out[18]), .IN3(
        divider_out[19]), .IN4(divider_out[1]), .Q(n535) );
  NOR4X0 U597 ( .IN1(n520), .IN2(n521), .IN3(n522), .IN4(n523), .QN(n519) );
  NOR4X0 U598 ( .IN1(n531), .IN2(n532), .IN3(n533), .IN4(n534), .QN(n530) );
  NAND4X0 U599 ( .IN1(divider_out[8]), .IN2(divider_out[3]), .IN3(
        divider_out[2]), .IN4(divider_out[1]), .QN(n527) );
  NAND2X1 U600 ( .IN1(n249), .IN2(n250), .QN(N435) );
  NAND2X1 U601 ( .IN1(n351), .IN2(n352), .QN(N384) );
  NAND2X1 U602 ( .IN1(n349), .IN2(n350), .QN(N385) );
  NAND2X1 U603 ( .IN1(n347), .IN2(n348), .QN(N386) );
  NAND2X1 U604 ( .IN1(n345), .IN2(n346), .QN(N387) );
  NAND2X1 U605 ( .IN1(n343), .IN2(n344), .QN(N388) );
  NAND2X1 U606 ( .IN1(n341), .IN2(n342), .QN(N389) );
  NAND2X1 U607 ( .IN1(n339), .IN2(n340), .QN(N390) );
  NAND2X1 U608 ( .IN1(n337), .IN2(n338), .QN(N391) );
  NAND2X1 U609 ( .IN1(n335), .IN2(n336), .QN(N392) );
  NAND2X1 U610 ( .IN1(n333), .IN2(n334), .QN(N393) );
  NAND2X1 U611 ( .IN1(n331), .IN2(n332), .QN(N394) );
  NAND2X1 U612 ( .IN1(n329), .IN2(n330), .QN(N395) );
  NAND2X1 U613 ( .IN1(n327), .IN2(n328), .QN(N396) );
  NAND2X1 U614 ( .IN1(n325), .IN2(n326), .QN(N397) );
  NAND2X1 U615 ( .IN1(n323), .IN2(n324), .QN(N398) );
  NAND2X1 U616 ( .IN1(n321), .IN2(n322), .QN(N399) );
  NAND2X1 U617 ( .IN1(n319), .IN2(n320), .QN(N400) );
  NAND2X1 U618 ( .IN1(n317), .IN2(n318), .QN(N401) );
  NAND2X1 U619 ( .IN1(n315), .IN2(n316), .QN(N402) );
  NAND2X1 U620 ( .IN1(n313), .IN2(n314), .QN(N403) );
  NAND2X1 U621 ( .IN1(n311), .IN2(n312), .QN(N404) );
  NAND2X1 U622 ( .IN1(n309), .IN2(n310), .QN(N405) );
  NAND2X1 U623 ( .IN1(n307), .IN2(n308), .QN(N406) );
  NAND2X1 U624 ( .IN1(n305), .IN2(n306), .QN(N407) );
  NAND2X1 U625 ( .IN1(n303), .IN2(n304), .QN(N408) );
  NAND2X1 U626 ( .IN1(n301), .IN2(n302), .QN(N409) );
  NAND2X1 U627 ( .IN1(n299), .IN2(n300), .QN(N410) );
  NAND2X1 U628 ( .IN1(n297), .IN2(n298), .QN(N411) );
  NAND2X1 U629 ( .IN1(n295), .IN2(n296), .QN(N412) );
  NAND2X1 U630 ( .IN1(n293), .IN2(n294), .QN(N413) );
  NAND2X1 U631 ( .IN1(n291), .IN2(n292), .QN(N414) );
  NAND2X1 U632 ( .IN1(n289), .IN2(n290), .QN(N415) );
  NAND2X1 U633 ( .IN1(n287), .IN2(n288), .QN(N416) );
  NAND2X1 U634 ( .IN1(n285), .IN2(n286), .QN(N417) );
  NAND2X1 U635 ( .IN1(n283), .IN2(n284), .QN(N418) );
  NAND2X1 U636 ( .IN1(n281), .IN2(n282), .QN(N419) );
  NAND2X1 U637 ( .IN1(n279), .IN2(n280), .QN(N420) );
  NAND2X1 U638 ( .IN1(n277), .IN2(n278), .QN(N421) );
  NAND2X1 U639 ( .IN1(n275), .IN2(n276), .QN(N422) );
  NAND2X1 U640 ( .IN1(n273), .IN2(n274), .QN(N423) );
  NAND2X1 U641 ( .IN1(n271), .IN2(n272), .QN(N424) );
  NAND2X1 U642 ( .IN1(n269), .IN2(n270), .QN(N425) );
  NAND2X1 U643 ( .IN1(n267), .IN2(n268), .QN(N426) );
  NAND2X1 U644 ( .IN1(n265), .IN2(n266), .QN(N427) );
  NAND2X1 U645 ( .IN1(n263), .IN2(n264), .QN(N428) );
  NAND2X1 U646 ( .IN1(n261), .IN2(n262), .QN(N429) );
  NAND2X1 U647 ( .IN1(n259), .IN2(n260), .QN(N430) );
  NAND2X1 U648 ( .IN1(n257), .IN2(n258), .QN(N431) );
  NAND2X1 U649 ( .IN1(n255), .IN2(n256), .QN(N432) );
  NAND2X1 U650 ( .IN1(n253), .IN2(n254), .QN(N433) );
  NAND2X1 U651 ( .IN1(n251), .IN2(n252), .QN(N434) );
  NAND2X1 U652 ( .IN1(n247), .IN2(n248), .QN(N436) );
  NAND2X1 U653 ( .IN1(n245), .IN2(n246), .QN(N437) );
  NAND2X1 U654 ( .IN1(n243), .IN2(n244), .QN(N438) );
  NAND2X1 U655 ( .IN1(n241), .IN2(n242), .QN(N439) );
  NAND2X1 U656 ( .IN1(n239), .IN2(n240), .QN(N440) );
  NAND2X1 U657 ( .IN1(n237), .IN2(n238), .QN(N441) );
  NAND2X1 U658 ( .IN1(n235), .IN2(n236), .QN(N442) );
  NAND2X1 U659 ( .IN1(n233), .IN2(n234), .QN(N443) );
  NAND2X1 U660 ( .IN1(n231), .IN2(n232), .QN(N444) );
  NAND2X1 U661 ( .IN1(n229), .IN2(n230), .QN(N445) );
  NAND2X1 U662 ( .IN1(n227), .IN2(n228), .QN(N446) );
  NAND2X1 U663 ( .IN1(data_tan[62]), .IN2(n649), .QN(n227) );
  NAND2X1 U664 ( .IN1(n225), .IN2(n226), .QN(N447) );
  INVX0 U665 ( .INP(n767), .ZN(n772) );
  INVX0 U666 ( .INP(n764), .ZN(n773) );
  NAND2X1 U667 ( .IN1(enable), .IN2(n819), .QN(n359) );
  INVX0 U668 ( .INP(rst), .ZN(n819) );
  INVX0 U669 ( .INP(degrees[20]), .ZN(n806) );
  INVX0 U670 ( .INP(degrees[23]), .ZN(n803) );
  INVX0 U671 ( .INP(degrees[21]), .ZN(n805) );
  INVX0 U672 ( .INP(degrees[17]), .ZN(n809) );
  INVX0 U673 ( .INP(degrees[1]), .ZN(n817) );
  INVX0 U674 ( .INP(degrees[18]), .ZN(n808) );
  INVX0 U675 ( .INP(degrees[0]), .ZN(n818) );
  INVX0 U676 ( .INP(degrees[12]), .ZN(n814) );
  INVX0 U677 ( .INP(degrees[10]), .ZN(n816) );
  INVX0 U678 ( .INP(degrees[24]), .ZN(n802) );
  INVX0 U679 ( .INP(degrees[27]), .ZN(n799) );
  INVX0 U680 ( .INP(degrees[25]), .ZN(n801) );
  INVX0 U681 ( .INP(degrees[13]), .ZN(n813) );
  INVX0 U682 ( .INP(degrees[16]), .ZN(n810) );
  INVX0 U683 ( .INP(degrees[14]), .ZN(n812) );
  INVX0 U684 ( .INP(degrees[7]), .ZN(n722) );
  INVX0 U685 ( .INP(actv[2]), .ZN(n822) );
  INVX0 U686 ( .INP(actv[1]), .ZN(n823) );
  INVX0 U687 ( .INP(actv[0]), .ZN(n824) );
  NOR4X0 U688 ( .IN1(n504), .IN2(n505), .IN3(n506), .IN4(n507), .QN(n498) );
  NOR4X0 U689 ( .IN1(n504), .IN2(n505), .IN3(n506), .IN4(n513), .QN(n509) );
  INVX0 U690 ( .INP(degrees[4]), .ZN(n770) );
  INVX0 U691 ( .INP(degrees[5]), .ZN(n771) );
  INVX0 U692 ( .INP(degrees[19]), .ZN(n807) );
  INVX0 U693 ( .INP(degrees[11]), .ZN(n815) );
  INVX0 U694 ( .INP(degrees[15]), .ZN(n811) );
  INVX0 U695 ( .INP(degrees[22]), .ZN(n804) );
  INVX0 U696 ( .INP(degrees[26]), .ZN(n800) );
  AO22X1 U697 ( .IN1(N194), .IN2(n678), .IN3(n639), .IN4(n679), .Q(n538) );
  INVX0 U698 ( .INP(divider_out[0]), .ZN(n796) );
  NAND2X0 U699 ( .IN1(n640), .IN2(n641), .QN(N355) );
  AOI221X1 U700 ( .IN1(divider_out[31]), .IN2(n663), .IN3(N157), .IN4(n672), 
        .IN5(n371), .QN(n640) );
  AOI221X1 U701 ( .IN1(n666), .IN2(degrees_tmp1[31]), .IN3(N258), .IN4(n670), 
        .IN5(n368), .QN(n641) );
  OR3X1 U702 ( .IN1(degrees_tmp1[14]), .IN2(degrees_tmp1[13]), .IN3(
        degrees_tmp1[12]), .Q(n685) );
  OA21X1 U703 ( .IN1(degrees_tmp1[5]), .IN2(degrees_tmp1[4]), .IN3(
        degrees_tmp1[6]), .Q(n683) );
  NAND2X0 U704 ( .IN1(degrees_tmp1[2]), .IN2(degrees_tmp1[3]), .QN(n681) );
  NAND4X0 U705 ( .IN1(n681), .IN2(n680), .IN3(n693), .IN4(n694), .QN(n682) );
  OA21X1 U706 ( .IN1(degrees_tmp1[7]), .IN2(n683), .IN3(n682), .Q(n684) );
  NOR4X0 U707 ( .IN1(n685), .IN2(n684), .IN3(degrees_tmp1[11]), .IN4(
        degrees_tmp1[10]), .QN(n692) );
  OR3X1 U708 ( .IN1(degrees_tmp1[20]), .IN2(degrees_tmp1[19]), .IN3(
        degrees_tmp1[18]), .Q(n686) );
  NOR4X0 U709 ( .IN1(n686), .IN2(degrees_tmp1[15]), .IN3(degrees_tmp1[17]), 
        .IN4(degrees_tmp1[16]), .QN(n691) );
  OR3X1 U710 ( .IN1(degrees_tmp1[26]), .IN2(degrees_tmp1[25]), .IN3(
        degrees_tmp1[24]), .Q(n687) );
  NOR4X0 U711 ( .IN1(n687), .IN2(degrees_tmp1[21]), .IN3(degrees_tmp1[23]), 
        .IN4(degrees_tmp1[22]), .QN(n690) );
  OR4X1 U712 ( .IN1(degrees_tmp1[31]), .IN2(degrees_tmp1[30]), .IN3(
        degrees_tmp1[9]), .IN4(degrees_tmp1[8]), .Q(n688) );
  NOR4X0 U713 ( .IN1(n688), .IN2(degrees_tmp1[27]), .IN3(degrees_tmp1[29]), 
        .IN4(degrees_tmp1[28]), .QN(n689) );
  NAND4X0 U714 ( .IN1(n692), .IN2(n691), .IN3(n690), .IN4(n689), .QN(N225) );
  OR3X1 U715 ( .IN1(divider_out[14]), .IN2(divider_out[13]), .IN3(
        divider_out[12]), .Q(n700) );
  OA21X1 U716 ( .IN1(divider_out[5]), .IN2(divider_out[4]), .IN3(
        divider_out[6]), .Q(n698) );
  NAND2X0 U717 ( .IN1(divider_out[2]), .IN2(divider_out[3]), .QN(n696) );
  NAND4X0 U718 ( .IN1(n696), .IN2(n695), .IN3(n739), .IN4(n708), .QN(n697) );
  OA21X1 U719 ( .IN1(divider_out[7]), .IN2(n698), .IN3(n697), .Q(n699) );
  NOR4X0 U720 ( .IN1(n700), .IN2(n699), .IN3(divider_out[11]), .IN4(
        divider_out[10]), .QN(n707) );
  OR3X1 U721 ( .IN1(divider_out[20]), .IN2(divider_out[19]), .IN3(
        divider_out[18]), .Q(n701) );
  NOR4X0 U722 ( .IN1(n701), .IN2(divider_out[15]), .IN3(divider_out[17]), 
        .IN4(divider_out[16]), .QN(n706) );
  OR3X1 U723 ( .IN1(divider_out[26]), .IN2(divider_out[25]), .IN3(
        divider_out[24]), .Q(n702) );
  NOR4X0 U724 ( .IN1(n702), .IN2(divider_out[21]), .IN3(divider_out[23]), 
        .IN4(divider_out[22]), .QN(n705) );
  OR4X1 U725 ( .IN1(divider_out[31]), .IN2(divider_out[30]), .IN3(
        divider_out[9]), .IN4(divider_out[8]), .Q(n703) );
  NOR4X0 U726 ( .IN1(n703), .IN2(divider_out[27]), .IN3(divider_out[29]), 
        .IN4(divider_out[28]), .QN(n704) );
  NAND4X0 U727 ( .IN1(n707), .IN2(n706), .IN3(n705), .IN4(n704), .QN(N54) );
  OR3X1 U728 ( .IN1(degrees[14]), .IN2(degrees[13]), .IN3(degrees[12]), .Q(
        n714) );
  OA21X1 U729 ( .IN1(degrees[5]), .IN2(degrees[4]), .IN3(degrees[6]), .Q(n712)
         );
  NAND2X0 U730 ( .IN1(degrees[2]), .IN2(degrees[3]), .QN(n710) );
  NAND3X0 U731 ( .IN1(degrees[1]), .IN2(degrees[0]), .IN3(degrees[3]), .QN(
        n709) );
  NAND4X0 U732 ( .IN1(n710), .IN2(n709), .IN3(n771), .IN4(n722), .QN(n711) );
  OA21X1 U733 ( .IN1(degrees[7]), .IN2(n712), .IN3(n711), .Q(n713) );
  NOR4X0 U734 ( .IN1(n714), .IN2(n713), .IN3(degrees[11]), .IN4(degrees[10]), 
        .QN(n721) );
  OR3X1 U735 ( .IN1(degrees[20]), .IN2(degrees[19]), .IN3(degrees[18]), .Q(
        n715) );
  NOR4X0 U736 ( .IN1(n715), .IN2(degrees[15]), .IN3(degrees[17]), .IN4(
        degrees[16]), .QN(n720) );
  OR3X1 U737 ( .IN1(degrees[26]), .IN2(degrees[25]), .IN3(degrees[24]), .Q(
        n716) );
  NOR4X0 U738 ( .IN1(n716), .IN2(degrees[21]), .IN3(degrees[23]), .IN4(
        degrees[22]), .QN(n719) );
  OR4X1 U739 ( .IN1(degrees[31]), .IN2(degrees[30]), .IN3(degrees[9]), .IN4(
        degrees[8]), .Q(n717) );
  NOR4X0 U740 ( .IN1(n717), .IN2(degrees[27]), .IN3(degrees[29]), .IN4(
        degrees[28]), .QN(n718) );
  NAND4X0 U741 ( .IN1(n721), .IN2(n720), .IN3(n719), .IN4(n718), .QN(N43) );
  NOR3X0 U742 ( .IN1(divider_out[31]), .IN2(divider_out[30]), .IN3(
        divider_out[29]), .QN(n731) );
  OR4X1 U743 ( .IN1(divider_out[14]), .IN2(divider_out[13]), .IN3(
        divider_out[9]), .IN4(divider_out[8]), .Q(n723) );
  NOR4X0 U744 ( .IN1(divider_out[12]), .IN2(divider_out[11]), .IN3(
        divider_out[10]), .IN4(n723), .QN(n730) );
  NOR2X0 U745 ( .IN1(divider_out[2]), .IN2(divider_out[3]), .QN(n733) );
  NOR3X0 U746 ( .IN1(divider_out[0]), .IN2(divider_out[3]), .IN3(
        divider_out[1]), .QN(n724) );
  NOR4X0 U747 ( .IN1(n733), .IN2(n724), .IN3(n738), .IN4(n739), .QN(n725) );
  NOR2X0 U748 ( .IN1(divider_out[6]), .IN2(n725), .QN(n727) );
  OR4X1 U749 ( .IN1(divider_out[19]), .IN2(divider_out[18]), .IN3(
        divider_out[21]), .IN4(divider_out[20]), .Q(n726) );
  NOR4X0 U750 ( .IN1(divider_out[17]), .IN2(divider_out[16]), .IN3(
        divider_out[15]), .IN4(n726), .QN(n735) );
  OA21X1 U751 ( .IN1(n727), .IN2(n708), .IN3(n735), .Q(n729) );
  OR4X1 U752 ( .IN1(divider_out[26]), .IN2(divider_out[25]), .IN3(
        divider_out[28]), .IN4(divider_out[27]), .Q(n728) );
  NOR4X0 U753 ( .IN1(divider_out[24]), .IN2(divider_out[23]), .IN3(
        divider_out[22]), .IN4(n728), .QN(n732) );
  NAND4X0 U754 ( .IN1(n731), .IN2(n730), .IN3(n729), .IN4(n732), .QN(N51) );
  NAND2X0 U755 ( .IN1(n731), .IN2(n730), .QN(n737) );
  NOR3X0 U756 ( .IN1(n739), .IN2(n733), .IN3(n738), .QN(n734) );
  OA21X1 U757 ( .IN1(n734), .IN2(divider_out[6]), .IN3(divider_out[7]), .Q(
        n736) );
  NOR4X0 U758 ( .IN1(n737), .IN2(n741), .IN3(n736), .IN4(n740), .QN(N55) );
  OR4X1 U759 ( .IN1(divider_out[5]), .IN2(divider_out[4]), .IN3(divider_out[7]), .IN4(divider_out[6]), .Q(n751) );
  AO21X1 U760 ( .IN1(divider_out[0]), .IN2(n752), .IN3(n751), .Q(n750) );
  OR2X1 U761 ( .IN1(divider_out[11]), .IN2(divider_out[10]), .Q(n742) );
  NOR4X0 U762 ( .IN1(n742), .IN2(divider_out[12]), .IN3(divider_out[14]), 
        .IN4(divider_out[13]), .QN(n749) );
  OR3X1 U763 ( .IN1(divider_out[20]), .IN2(divider_out[19]), .IN3(
        divider_out[18]), .Q(n743) );
  NOR4X0 U764 ( .IN1(n743), .IN2(divider_out[15]), .IN3(divider_out[17]), 
        .IN4(divider_out[16]), .QN(n748) );
  OR3X1 U765 ( .IN1(divider_out[26]), .IN2(divider_out[25]), .IN3(
        divider_out[24]), .Q(n744) );
  NOR4X0 U766 ( .IN1(n744), .IN2(divider_out[21]), .IN3(divider_out[23]), 
        .IN4(divider_out[22]), .QN(n747) );
  OR3X1 U767 ( .IN1(divider_out[9]), .IN2(divider_out[31]), .IN3(
        divider_out[30]), .Q(n745) );
  NOR4X0 U768 ( .IN1(n745), .IN2(divider_out[27]), .IN3(divider_out[29]), 
        .IN4(divider_out[28]), .QN(n746) );
  NAND4X0 U769 ( .IN1(n749), .IN2(n748), .IN3(n747), .IN4(n746), .QN(n753) );
  AO21X1 U770 ( .IN1(divider_out[8]), .IN2(n750), .IN3(n753), .Q(N50) );
  OA21X1 U771 ( .IN1(n752), .IN2(n751), .IN3(divider_out[8]), .Q(n754) );
  NOR2X0 U772 ( .IN1(n754), .IN2(n753), .QN(N52) );
  NOR3X0 U773 ( .IN1(degrees[31]), .IN2(degrees[30]), .IN3(degrees[29]), .QN(
        n763) );
  OR4X1 U774 ( .IN1(degrees[14]), .IN2(degrees[13]), .IN3(degrees[9]), .IN4(
        degrees[8]), .Q(n755) );
  NOR4X0 U775 ( .IN1(degrees[12]), .IN2(degrees[11]), .IN3(degrees[10]), .IN4(
        n755), .QN(n762) );
  NOR2X0 U776 ( .IN1(degrees[2]), .IN2(degrees[3]), .QN(n765) );
  NOR3X0 U777 ( .IN1(degrees[0]), .IN2(degrees[3]), .IN3(degrees[1]), .QN(n756) );
  NOR4X0 U778 ( .IN1(n765), .IN2(n756), .IN3(n770), .IN4(n771), .QN(n757) );
  NOR2X0 U779 ( .IN1(degrees[6]), .IN2(n757), .QN(n759) );
  OR4X1 U780 ( .IN1(degrees[19]), .IN2(degrees[18]), .IN3(degrees[21]), .IN4(
        degrees[20]), .Q(n758) );
  NOR4X0 U781 ( .IN1(degrees[17]), .IN2(degrees[16]), .IN3(degrees[15]), .IN4(
        n758), .QN(n767) );
  OA21X1 U782 ( .IN1(n759), .IN2(n722), .IN3(n767), .Q(n761) );
  OR4X1 U783 ( .IN1(degrees[26]), .IN2(degrees[25]), .IN3(degrees[28]), .IN4(
        degrees[27]), .Q(n760) );
  NOR4X0 U784 ( .IN1(degrees[24]), .IN2(degrees[23]), .IN3(degrees[22]), .IN4(
        n760), .QN(n764) );
  NAND4X0 U785 ( .IN1(n763), .IN2(n762), .IN3(n761), .IN4(n764), .QN(N40) );
  NAND2X0 U786 ( .IN1(n763), .IN2(n762), .QN(n769) );
  NOR3X0 U787 ( .IN1(n771), .IN2(n765), .IN3(n770), .QN(n766) );
  OA21X1 U788 ( .IN1(n766), .IN2(degrees[6]), .IN3(degrees[7]), .Q(n768) );
  NOR4X0 U789 ( .IN1(n769), .IN2(n773), .IN3(n768), .IN4(n772), .QN(N44) );
  OR2X1 U790 ( .IN1(degrees[3]), .IN2(degrees[4]), .Q(n774) );
  AND4X1 U791 ( .IN1(degrees[6]), .IN2(degrees[5]), .IN3(degrees[8]), .IN4(
        n774), .Q(n786) );
  OR4X1 U792 ( .IN1(degrees[1]), .IN2(degrees[0]), .IN3(degrees[4]), .IN4(
        degrees[2]), .Q(n784) );
  OR3X1 U793 ( .IN1(degrees[14]), .IN2(degrees[13]), .IN3(degrees[12]), .Q(
        n776) );
  AND2X1 U794 ( .IN1(degrees[8]), .IN2(degrees[7]), .Q(n775) );
  NOR4X0 U795 ( .IN1(n776), .IN2(n775), .IN3(degrees[11]), .IN4(degrees[10]), 
        .QN(n783) );
  OR3X1 U796 ( .IN1(degrees[20]), .IN2(degrees[19]), .IN3(degrees[18]), .Q(
        n777) );
  NOR4X0 U797 ( .IN1(n777), .IN2(degrees[15]), .IN3(degrees[17]), .IN4(
        degrees[16]), .QN(n782) );
  OR3X1 U798 ( .IN1(degrees[26]), .IN2(degrees[25]), .IN3(degrees[24]), .Q(
        n778) );
  NOR4X0 U799 ( .IN1(n778), .IN2(degrees[21]), .IN3(degrees[23]), .IN4(
        degrees[22]), .QN(n781) );
  OR3X1 U800 ( .IN1(degrees[9]), .IN2(degrees[31]), .IN3(degrees[30]), .Q(n779) );
  NOR4X0 U801 ( .IN1(n779), .IN2(degrees[27]), .IN3(degrees[29]), .IN4(
        degrees[28]), .QN(n780) );
  NAND4X0 U802 ( .IN1(n783), .IN2(n782), .IN3(n781), .IN4(n780), .QN(n785) );
  AO21X1 U803 ( .IN1(n786), .IN2(n784), .IN3(n785), .Q(N39) );
  NOR2X0 U804 ( .IN1(n786), .IN2(n785), .QN(N41) );
endmodule

